module Memory(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_1(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_2(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_3(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_4(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_5(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_6(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_7(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_8(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_8.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_9(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_9.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_10(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_10.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_11(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_11.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_12(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_12.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_13(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_13.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_14(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_14.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_15(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_15.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_16(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_16.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_17(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_17.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_18(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_18.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_19(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_19.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_20(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_20.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_21(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_21.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_22(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_22.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_23(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_23.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_24(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_24.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_25(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_25.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_26(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_26.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_27(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_27.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_28(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_28.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_29(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_29.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_30(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_30.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_31(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_31.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_64(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead,
  input         io_writeEnable,
  input  [4:0]  io_dataWrite
);
  wire  RamSpWf_clk; // @[Memory.scala 57:26]
  wire  RamSpWf_we; // @[Memory.scala 57:26]
  wire  RamSpWf_en; // @[Memory.scala 57:26]
  wire [10:0] RamSpWf_addr; // @[Memory.scala 57:26]
  wire [4:0] RamSpWf_di; // @[Memory.scala 57:26]
  wire [4:0] RamSpWf_dout; // @[Memory.scala 57:26]
  RamSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5)) RamSpWf ( // @[Memory.scala 57:26]
    .clk(RamSpWf_clk),
    .we(RamSpWf_we),
    .en(RamSpWf_en),
    .addr(RamSpWf_addr),
    .di(RamSpWf_di),
    .dout(RamSpWf_dout)
  );
  assign io_dataRead = RamSpWf_dout; // @[Memory.scala 63:17]
  assign RamSpWf_clk = clock; // @[Memory.scala 58:21]
  assign RamSpWf_we = io_writeEnable; // @[Memory.scala 59:20]
  assign RamSpWf_en = 1'h1; // @[Memory.scala 60:20]
  assign RamSpWf_addr = io_address; // @[Memory.scala 61:22]
  assign RamSpWf_di = io_dataWrite; // @[Memory.scala 62:20]
endmodule
module Memory_68(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [10:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5), .LOAD_FILE("memory_init/backbuffer_init0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 5'h0; // @[Memory.scala 70:20]
endmodule
module Memory_69(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [10:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5), .LOAD_FILE("memory_init/backbuffer_init1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 5'h0; // @[Memory.scala 70:20]
endmodule
module Memory_70(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_71(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_72(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_73(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_74(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_75(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_76(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_77(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_78(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_8.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_79(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_9.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_80(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_10.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_81(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_11.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_82(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_12.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_83(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_13.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_84(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_14.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_85(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_15.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_86(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_16.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_87(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_17.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_88(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_18.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_89(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_19.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_90(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_20.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_91(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_21.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_92(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_22.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_93(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_23.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_94(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_24.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_95(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_25.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_96(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_26.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_97(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_27.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_98(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_28.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_99(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_29.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_100(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_30.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_101(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_31.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_102(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_32.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_103(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_33.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_104(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_34.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_105(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_35.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_106(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_36.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_107(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_37.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_108(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_38.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_109(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_39.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_110(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_40.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_111(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_41.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_112(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_42.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_113(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_43.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_114(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_44.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_115(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_45.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_116(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_46.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_117(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_47.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_118(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_48.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_119(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_49.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_120(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_50.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_121(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_51.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_122(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_52.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_123(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_53.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_124(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_54.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_125(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_55.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_126(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_56.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_127(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_57.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_128(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_58.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_129(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_59.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_130(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_60.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_131(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_61.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_132(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_62.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_133(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_63.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_134(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_64.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_135(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_65.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_136(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_66.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_137(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_67.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_138(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_68.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_139(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_69.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_140(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_70.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_141(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_71.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_142(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_72.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_143(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_73.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_144(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_74.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_145(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_75.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_146(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_76.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_147(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_77.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_148(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_78.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_149(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_79.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_150(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_80.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_151(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_81.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_152(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_82.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_153(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_83.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_154(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_84.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_155(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_85.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_156(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_86.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_157(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_87.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_158(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_88.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_159(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_89.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_160(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_90.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_161(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_91.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_162(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_92.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_163(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_93.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_164(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_94.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_165(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_95.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_166(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_96.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_167(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_97.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_168(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_98.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_169(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_99.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_170(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_100.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_171(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_101.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_172(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_102.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_173(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_103.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_174(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_104.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_175(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_105.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_176(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_106.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_177(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_107.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_178(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_108.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_179(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_109.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_180(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_110.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_181(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_111.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_182(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_112.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_183(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_113.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_184(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_114.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_185(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_115.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_186(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_116.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_187(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_117.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_188(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_118.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_189(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_119.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_190(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_120.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_191(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_121.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_192(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_122.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_193(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_123.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_194(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_124.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_195(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_125.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_196(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_126.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_197(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_127.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_198(
  input         clock,
  input  [11:0] io_address
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [11:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [14:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [14:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(12), .DATA_WIDTH(15), .LOAD_FILE("memory_init/rotation45deg.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 15'h0; // @[Memory.scala 70:20]
endmodule
module MultiHotPriortyReductionTree(
  input  [6:0] io_dataInput_0,
  input  [6:0] io_dataInput_1,
  input  [6:0] io_dataInput_2,
  input  [6:0] io_dataInput_3,
  input  [6:0] io_dataInput_4,
  input  [6:0] io_dataInput_5,
  input  [6:0] io_dataInput_6,
  input  [6:0] io_dataInput_7,
  input  [6:0] io_dataInput_8,
  input  [6:0] io_dataInput_9,
  input  [6:0] io_dataInput_10,
  input  [6:0] io_dataInput_11,
  input  [6:0] io_dataInput_12,
  input  [6:0] io_dataInput_13,
  input  [6:0] io_dataInput_14,
  input  [6:0] io_dataInput_15,
  input  [6:0] io_dataInput_16,
  input  [6:0] io_dataInput_17,
  input  [6:0] io_dataInput_18,
  input  [6:0] io_dataInput_19,
  input  [6:0] io_dataInput_20,
  input  [6:0] io_dataInput_21,
  input  [6:0] io_dataInput_22,
  input  [6:0] io_dataInput_23,
  input  [6:0] io_dataInput_24,
  input  [6:0] io_dataInput_25,
  input  [6:0] io_dataInput_26,
  input  [6:0] io_dataInput_27,
  input  [6:0] io_dataInput_28,
  input  [6:0] io_dataInput_29,
  input  [6:0] io_dataInput_30,
  input  [6:0] io_dataInput_31,
  input  [6:0] io_dataInput_32,
  input  [6:0] io_dataInput_33,
  input  [6:0] io_dataInput_34,
  input  [6:0] io_dataInput_35,
  input  [6:0] io_dataInput_36,
  input  [6:0] io_dataInput_37,
  input  [6:0] io_dataInput_38,
  input  [6:0] io_dataInput_39,
  input  [6:0] io_dataInput_40,
  input  [6:0] io_dataInput_41,
  input  [6:0] io_dataInput_42,
  input  [6:0] io_dataInput_43,
  input  [6:0] io_dataInput_44,
  input  [6:0] io_dataInput_45,
  input  [6:0] io_dataInput_46,
  input  [6:0] io_dataInput_47,
  input  [6:0] io_dataInput_48,
  input  [6:0] io_dataInput_49,
  input  [6:0] io_dataInput_50,
  input  [6:0] io_dataInput_51,
  input  [6:0] io_dataInput_52,
  input  [6:0] io_dataInput_53,
  input  [6:0] io_dataInput_54,
  input  [6:0] io_dataInput_55,
  input  [6:0] io_dataInput_56,
  input  [6:0] io_dataInput_57,
  input  [6:0] io_dataInput_58,
  input  [6:0] io_dataInput_59,
  input  [6:0] io_dataInput_60,
  input  [6:0] io_dataInput_61,
  input  [6:0] io_dataInput_62,
  input  [6:0] io_dataInput_63,
  input  [6:0] io_dataInput_64,
  input  [6:0] io_dataInput_65,
  input  [6:0] io_dataInput_66,
  input  [6:0] io_dataInput_67,
  input  [6:0] io_dataInput_68,
  input  [6:0] io_dataInput_69,
  input  [6:0] io_dataInput_70,
  input  [6:0] io_dataInput_71,
  input  [6:0] io_dataInput_72,
  input  [6:0] io_dataInput_73,
  input  [6:0] io_dataInput_74,
  input  [6:0] io_dataInput_75,
  input  [6:0] io_dataInput_76,
  input  [6:0] io_dataInput_77,
  input  [6:0] io_dataInput_78,
  input  [6:0] io_dataInput_79,
  input  [6:0] io_dataInput_80,
  input  [6:0] io_dataInput_81,
  input  [6:0] io_dataInput_82,
  input  [6:0] io_dataInput_83,
  input  [6:0] io_dataInput_84,
  input  [6:0] io_dataInput_85,
  input  [6:0] io_dataInput_86,
  input  [6:0] io_dataInput_87,
  input  [6:0] io_dataInput_88,
  input  [6:0] io_dataInput_89,
  input  [6:0] io_dataInput_90,
  input  [6:0] io_dataInput_91,
  input  [6:0] io_dataInput_92,
  input  [6:0] io_dataInput_93,
  input  [6:0] io_dataInput_94,
  input  [6:0] io_dataInput_95,
  input  [6:0] io_dataInput_96,
  input  [6:0] io_dataInput_97,
  input  [6:0] io_dataInput_98,
  input  [6:0] io_dataInput_99,
  input  [6:0] io_dataInput_100,
  input  [6:0] io_dataInput_101,
  input  [6:0] io_dataInput_102,
  input  [6:0] io_dataInput_103,
  input  [6:0] io_dataInput_104,
  input  [6:0] io_dataInput_105,
  input  [6:0] io_dataInput_106,
  input  [6:0] io_dataInput_107,
  input  [6:0] io_dataInput_108,
  input  [6:0] io_dataInput_109,
  input  [6:0] io_dataInput_110,
  input  [6:0] io_dataInput_111,
  input  [6:0] io_dataInput_112,
  input  [6:0] io_dataInput_113,
  input  [6:0] io_dataInput_114,
  input  [6:0] io_dataInput_115,
  input  [6:0] io_dataInput_116,
  input  [6:0] io_dataInput_117,
  input  [6:0] io_dataInput_118,
  input  [6:0] io_dataInput_119,
  input  [6:0] io_dataInput_120,
  input  [6:0] io_dataInput_121,
  input  [6:0] io_dataInput_122,
  input  [6:0] io_dataInput_123,
  input  [6:0] io_dataInput_124,
  input  [6:0] io_dataInput_125,
  input  [6:0] io_dataInput_126,
  input  [6:0] io_dataInput_127,
  input        io_selectInput_0,
  input        io_selectInput_1,
  input        io_selectInput_2,
  input        io_selectInput_3,
  input        io_selectInput_4,
  input        io_selectInput_5,
  input        io_selectInput_6,
  input        io_selectInput_7,
  input        io_selectInput_8,
  input        io_selectInput_9,
  input        io_selectInput_10,
  input        io_selectInput_11,
  input        io_selectInput_12,
  input        io_selectInput_13,
  input        io_selectInput_14,
  input        io_selectInput_15,
  input        io_selectInput_16,
  input        io_selectInput_17,
  input        io_selectInput_18,
  input        io_selectInput_19,
  input        io_selectInput_20,
  input        io_selectInput_21,
  input        io_selectInput_22,
  input        io_selectInput_23,
  input        io_selectInput_24,
  input        io_selectInput_25,
  input        io_selectInput_26,
  input        io_selectInput_27,
  input        io_selectInput_28,
  input        io_selectInput_29,
  input        io_selectInput_30,
  input        io_selectInput_31,
  input        io_selectInput_32,
  input        io_selectInput_33,
  input        io_selectInput_34,
  input        io_selectInput_35,
  input        io_selectInput_36,
  input        io_selectInput_37,
  input        io_selectInput_38,
  input        io_selectInput_39,
  input        io_selectInput_40,
  input        io_selectInput_41,
  input        io_selectInput_42,
  input        io_selectInput_43,
  input        io_selectInput_44,
  input        io_selectInput_45,
  input        io_selectInput_46,
  input        io_selectInput_47,
  input        io_selectInput_48,
  input        io_selectInput_49,
  input        io_selectInput_50,
  input        io_selectInput_51,
  input        io_selectInput_52,
  input        io_selectInput_53,
  input        io_selectInput_54,
  input        io_selectInput_55,
  input        io_selectInput_56,
  input        io_selectInput_57,
  input        io_selectInput_58,
  input        io_selectInput_59,
  input        io_selectInput_60,
  input        io_selectInput_61,
  input        io_selectInput_62,
  input        io_selectInput_63,
  input        io_selectInput_64,
  input        io_selectInput_65,
  input        io_selectInput_66,
  input        io_selectInput_67,
  input        io_selectInput_68,
  input        io_selectInput_69,
  input        io_selectInput_70,
  input        io_selectInput_71,
  input        io_selectInput_72,
  input        io_selectInput_73,
  input        io_selectInput_74,
  input        io_selectInput_75,
  input        io_selectInput_76,
  input        io_selectInput_77,
  input        io_selectInput_78,
  input        io_selectInput_79,
  input        io_selectInput_80,
  input        io_selectInput_81,
  input        io_selectInput_82,
  input        io_selectInput_83,
  input        io_selectInput_84,
  input        io_selectInput_85,
  input        io_selectInput_86,
  input        io_selectInput_87,
  input        io_selectInput_88,
  input        io_selectInput_89,
  input        io_selectInput_90,
  input        io_selectInput_91,
  input        io_selectInput_92,
  input        io_selectInput_93,
  input        io_selectInput_94,
  input        io_selectInput_95,
  input        io_selectInput_96,
  input        io_selectInput_97,
  input        io_selectInput_98,
  input        io_selectInput_99,
  input        io_selectInput_100,
  input        io_selectInput_101,
  input        io_selectInput_102,
  input        io_selectInput_103,
  input        io_selectInput_104,
  input        io_selectInput_105,
  input        io_selectInput_106,
  input        io_selectInput_107,
  input        io_selectInput_108,
  input        io_selectInput_109,
  input        io_selectInput_110,
  input        io_selectInput_111,
  input        io_selectInput_112,
  input        io_selectInput_113,
  input        io_selectInput_114,
  input        io_selectInput_115,
  input        io_selectInput_116,
  input        io_selectInput_117,
  input        io_selectInput_118,
  input        io_selectInput_119,
  input        io_selectInput_120,
  input        io_selectInput_121,
  input        io_selectInput_122,
  input        io_selectInput_123,
  input        io_selectInput_124,
  input        io_selectInput_125,
  input        io_selectInput_126,
  input        io_selectInput_127,
  output [6:0] io_dataOutput,
  output       io_selectOutput,
  output [6:0] io_indexOutput
);
  wire  selectNodeOutputs_63 = io_selectInput_0 | io_selectInput_1; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_64 = io_selectInput_2 | io_selectInput_3; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_31 = selectNodeOutputs_63 | selectNodeOutputs_64; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_65 = io_selectInput_4 | io_selectInput_5; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_66 = io_selectInput_6 | io_selectInput_7; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_32 = selectNodeOutputs_65 | selectNodeOutputs_66; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_15 = selectNodeOutputs_31 | selectNodeOutputs_32; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_67 = io_selectInput_8 | io_selectInput_9; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_68 = io_selectInput_10 | io_selectInput_11; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_33 = selectNodeOutputs_67 | selectNodeOutputs_68; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_69 = io_selectInput_12 | io_selectInput_13; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_70 = io_selectInput_14 | io_selectInput_15; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_34 = selectNodeOutputs_69 | selectNodeOutputs_70; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_16 = selectNodeOutputs_33 | selectNodeOutputs_34; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_7 = selectNodeOutputs_15 | selectNodeOutputs_16; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_71 = io_selectInput_16 | io_selectInput_17; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_72 = io_selectInput_18 | io_selectInput_19; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_35 = selectNodeOutputs_71 | selectNodeOutputs_72; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_73 = io_selectInput_20 | io_selectInput_21; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_74 = io_selectInput_22 | io_selectInput_23; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_36 = selectNodeOutputs_73 | selectNodeOutputs_74; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_17 = selectNodeOutputs_35 | selectNodeOutputs_36; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_75 = io_selectInput_24 | io_selectInput_25; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_76 = io_selectInput_26 | io_selectInput_27; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_37 = selectNodeOutputs_75 | selectNodeOutputs_76; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_77 = io_selectInput_28 | io_selectInput_29; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_78 = io_selectInput_30 | io_selectInput_31; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_38 = selectNodeOutputs_77 | selectNodeOutputs_78; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_18 = selectNodeOutputs_37 | selectNodeOutputs_38; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_8 = selectNodeOutputs_17 | selectNodeOutputs_18; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_3 = selectNodeOutputs_7 | selectNodeOutputs_8; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_79 = io_selectInput_32 | io_selectInput_33; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_80 = io_selectInput_34 | io_selectInput_35; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_39 = selectNodeOutputs_79 | selectNodeOutputs_80; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_81 = io_selectInput_36 | io_selectInput_37; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_82 = io_selectInput_38 | io_selectInput_39; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_40 = selectNodeOutputs_81 | selectNodeOutputs_82; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_19 = selectNodeOutputs_39 | selectNodeOutputs_40; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_83 = io_selectInput_40 | io_selectInput_41; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_84 = io_selectInput_42 | io_selectInput_43; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_41 = selectNodeOutputs_83 | selectNodeOutputs_84; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_85 = io_selectInput_44 | io_selectInput_45; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_86 = io_selectInput_46 | io_selectInput_47; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_42 = selectNodeOutputs_85 | selectNodeOutputs_86; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_20 = selectNodeOutputs_41 | selectNodeOutputs_42; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_9 = selectNodeOutputs_19 | selectNodeOutputs_20; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_87 = io_selectInput_48 | io_selectInput_49; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_88 = io_selectInput_50 | io_selectInput_51; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_43 = selectNodeOutputs_87 | selectNodeOutputs_88; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_89 = io_selectInput_52 | io_selectInput_53; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_90 = io_selectInput_54 | io_selectInput_55; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_44 = selectNodeOutputs_89 | selectNodeOutputs_90; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_21 = selectNodeOutputs_43 | selectNodeOutputs_44; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_91 = io_selectInput_56 | io_selectInput_57; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_92 = io_selectInput_58 | io_selectInput_59; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_45 = selectNodeOutputs_91 | selectNodeOutputs_92; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_93 = io_selectInput_60 | io_selectInput_61; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_94 = io_selectInput_62 | io_selectInput_63; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_46 = selectNodeOutputs_93 | selectNodeOutputs_94; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_22 = selectNodeOutputs_45 | selectNodeOutputs_46; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_10 = selectNodeOutputs_21 | selectNodeOutputs_22; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_4 = selectNodeOutputs_9 | selectNodeOutputs_10; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_1 = selectNodeOutputs_3 | selectNodeOutputs_4; // @[GameUtilities.scala 92:54]
  wire [6:0] dataNodeOutputs_63 = io_selectInput_0 ? io_dataInput_0 : io_dataInput_1; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_64 = io_selectInput_2 ? io_dataInput_2 : io_dataInput_3; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_31 = selectNodeOutputs_63 ? dataNodeOutputs_63 : dataNodeOutputs_64; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_65 = io_selectInput_4 ? io_dataInput_4 : io_dataInput_5; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_66 = io_selectInput_6 ? io_dataInput_6 : io_dataInput_7; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_32 = selectNodeOutputs_65 ? dataNodeOutputs_65 : dataNodeOutputs_66; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_15 = selectNodeOutputs_31 ? dataNodeOutputs_31 : dataNodeOutputs_32; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_67 = io_selectInput_8 ? io_dataInput_8 : io_dataInput_9; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_68 = io_selectInput_10 ? io_dataInput_10 : io_dataInput_11; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_33 = selectNodeOutputs_67 ? dataNodeOutputs_67 : dataNodeOutputs_68; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_69 = io_selectInput_12 ? io_dataInput_12 : io_dataInput_13; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_70 = io_selectInput_14 ? io_dataInput_14 : io_dataInput_15; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_34 = selectNodeOutputs_69 ? dataNodeOutputs_69 : dataNodeOutputs_70; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_16 = selectNodeOutputs_33 ? dataNodeOutputs_33 : dataNodeOutputs_34; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_7 = selectNodeOutputs_15 ? dataNodeOutputs_15 : dataNodeOutputs_16; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_71 = io_selectInput_16 ? io_dataInput_16 : io_dataInput_17; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_72 = io_selectInput_18 ? io_dataInput_18 : io_dataInput_19; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_35 = selectNodeOutputs_71 ? dataNodeOutputs_71 : dataNodeOutputs_72; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_73 = io_selectInput_20 ? io_dataInput_20 : io_dataInput_21; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_74 = io_selectInput_22 ? io_dataInput_22 : io_dataInput_23; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_36 = selectNodeOutputs_73 ? dataNodeOutputs_73 : dataNodeOutputs_74; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_17 = selectNodeOutputs_35 ? dataNodeOutputs_35 : dataNodeOutputs_36; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_75 = io_selectInput_24 ? io_dataInput_24 : io_dataInput_25; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_76 = io_selectInput_26 ? io_dataInput_26 : io_dataInput_27; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_37 = selectNodeOutputs_75 ? dataNodeOutputs_75 : dataNodeOutputs_76; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_77 = io_selectInput_28 ? io_dataInput_28 : io_dataInput_29; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_78 = io_selectInput_30 ? io_dataInput_30 : io_dataInput_31; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_38 = selectNodeOutputs_77 ? dataNodeOutputs_77 : dataNodeOutputs_78; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_18 = selectNodeOutputs_37 ? dataNodeOutputs_37 : dataNodeOutputs_38; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_8 = selectNodeOutputs_17 ? dataNodeOutputs_17 : dataNodeOutputs_18; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_3 = selectNodeOutputs_7 ? dataNodeOutputs_7 : dataNodeOutputs_8; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_79 = io_selectInput_32 ? io_dataInput_32 : io_dataInput_33; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_80 = io_selectInput_34 ? io_dataInput_34 : io_dataInput_35; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_39 = selectNodeOutputs_79 ? dataNodeOutputs_79 : dataNodeOutputs_80; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_81 = io_selectInput_36 ? io_dataInput_36 : io_dataInput_37; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_82 = io_selectInput_38 ? io_dataInput_38 : io_dataInput_39; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_40 = selectNodeOutputs_81 ? dataNodeOutputs_81 : dataNodeOutputs_82; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_19 = selectNodeOutputs_39 ? dataNodeOutputs_39 : dataNodeOutputs_40; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_83 = io_selectInput_40 ? io_dataInput_40 : io_dataInput_41; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_84 = io_selectInput_42 ? io_dataInput_42 : io_dataInput_43; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_41 = selectNodeOutputs_83 ? dataNodeOutputs_83 : dataNodeOutputs_84; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_85 = io_selectInput_44 ? io_dataInput_44 : io_dataInput_45; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_86 = io_selectInput_46 ? io_dataInput_46 : io_dataInput_47; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_42 = selectNodeOutputs_85 ? dataNodeOutputs_85 : dataNodeOutputs_86; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_20 = selectNodeOutputs_41 ? dataNodeOutputs_41 : dataNodeOutputs_42; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_9 = selectNodeOutputs_19 ? dataNodeOutputs_19 : dataNodeOutputs_20; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_87 = io_selectInput_48 ? io_dataInput_48 : io_dataInput_49; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_88 = io_selectInput_50 ? io_dataInput_50 : io_dataInput_51; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_43 = selectNodeOutputs_87 ? dataNodeOutputs_87 : dataNodeOutputs_88; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_89 = io_selectInput_52 ? io_dataInput_52 : io_dataInput_53; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_90 = io_selectInput_54 ? io_dataInput_54 : io_dataInput_55; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_44 = selectNodeOutputs_89 ? dataNodeOutputs_89 : dataNodeOutputs_90; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_21 = selectNodeOutputs_43 ? dataNodeOutputs_43 : dataNodeOutputs_44; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_91 = io_selectInput_56 ? io_dataInput_56 : io_dataInput_57; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_92 = io_selectInput_58 ? io_dataInput_58 : io_dataInput_59; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_45 = selectNodeOutputs_91 ? dataNodeOutputs_91 : dataNodeOutputs_92; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_93 = io_selectInput_60 ? io_dataInput_60 : io_dataInput_61; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_94 = io_selectInput_62 ? io_dataInput_62 : io_dataInput_63; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_46 = selectNodeOutputs_93 ? dataNodeOutputs_93 : dataNodeOutputs_94; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_22 = selectNodeOutputs_45 ? dataNodeOutputs_45 : dataNodeOutputs_46; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_10 = selectNodeOutputs_21 ? dataNodeOutputs_21 : dataNodeOutputs_22; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_4 = selectNodeOutputs_9 ? dataNodeOutputs_9 : dataNodeOutputs_10; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_1 = selectNodeOutputs_3 ? dataNodeOutputs_3 : dataNodeOutputs_4; // @[GameUtilities.scala 91:34]
  wire  selectNodeOutputs_95 = io_selectInput_64 | io_selectInput_65; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_96 = io_selectInput_66 | io_selectInput_67; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_47 = selectNodeOutputs_95 | selectNodeOutputs_96; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_97 = io_selectInput_68 | io_selectInput_69; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_98 = io_selectInput_70 | io_selectInput_71; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_48 = selectNodeOutputs_97 | selectNodeOutputs_98; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_23 = selectNodeOutputs_47 | selectNodeOutputs_48; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_99 = io_selectInput_72 | io_selectInput_73; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_100 = io_selectInput_74 | io_selectInput_75; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_49 = selectNodeOutputs_99 | selectNodeOutputs_100; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_101 = io_selectInput_76 | io_selectInput_77; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_102 = io_selectInput_78 | io_selectInput_79; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_50 = selectNodeOutputs_101 | selectNodeOutputs_102; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_24 = selectNodeOutputs_49 | selectNodeOutputs_50; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_11 = selectNodeOutputs_23 | selectNodeOutputs_24; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_103 = io_selectInput_80 | io_selectInput_81; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_104 = io_selectInput_82 | io_selectInput_83; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_51 = selectNodeOutputs_103 | selectNodeOutputs_104; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_105 = io_selectInput_84 | io_selectInput_85; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_106 = io_selectInput_86 | io_selectInput_87; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_52 = selectNodeOutputs_105 | selectNodeOutputs_106; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_25 = selectNodeOutputs_51 | selectNodeOutputs_52; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_107 = io_selectInput_88 | io_selectInput_89; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_108 = io_selectInput_90 | io_selectInput_91; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_53 = selectNodeOutputs_107 | selectNodeOutputs_108; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_109 = io_selectInput_92 | io_selectInput_93; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_110 = io_selectInput_94 | io_selectInput_95; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_54 = selectNodeOutputs_109 | selectNodeOutputs_110; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_26 = selectNodeOutputs_53 | selectNodeOutputs_54; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_12 = selectNodeOutputs_25 | selectNodeOutputs_26; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_5 = selectNodeOutputs_11 | selectNodeOutputs_12; // @[GameUtilities.scala 92:54]
  wire [6:0] dataNodeOutputs_95 = io_selectInput_64 ? io_dataInput_64 : io_dataInput_65; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_96 = io_selectInput_66 ? io_dataInput_66 : io_dataInput_67; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_47 = selectNodeOutputs_95 ? dataNodeOutputs_95 : dataNodeOutputs_96; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_97 = io_selectInput_68 ? io_dataInput_68 : io_dataInput_69; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_98 = io_selectInput_70 ? io_dataInput_70 : io_dataInput_71; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_48 = selectNodeOutputs_97 ? dataNodeOutputs_97 : dataNodeOutputs_98; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_23 = selectNodeOutputs_47 ? dataNodeOutputs_47 : dataNodeOutputs_48; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_99 = io_selectInput_72 ? io_dataInput_72 : io_dataInput_73; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_100 = io_selectInput_74 ? io_dataInput_74 : io_dataInput_75; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_49 = selectNodeOutputs_99 ? dataNodeOutputs_99 : dataNodeOutputs_100; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_101 = io_selectInput_76 ? io_dataInput_76 : io_dataInput_77; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_102 = io_selectInput_78 ? io_dataInput_78 : io_dataInput_79; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_50 = selectNodeOutputs_101 ? dataNodeOutputs_101 : dataNodeOutputs_102; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_24 = selectNodeOutputs_49 ? dataNodeOutputs_49 : dataNodeOutputs_50; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_11 = selectNodeOutputs_23 ? dataNodeOutputs_23 : dataNodeOutputs_24; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_103 = io_selectInput_80 ? io_dataInput_80 : io_dataInput_81; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_104 = io_selectInput_82 ? io_dataInput_82 : io_dataInput_83; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_51 = selectNodeOutputs_103 ? dataNodeOutputs_103 : dataNodeOutputs_104; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_105 = io_selectInput_84 ? io_dataInput_84 : io_dataInput_85; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_106 = io_selectInput_86 ? io_dataInput_86 : io_dataInput_87; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_52 = selectNodeOutputs_105 ? dataNodeOutputs_105 : dataNodeOutputs_106; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_25 = selectNodeOutputs_51 ? dataNodeOutputs_51 : dataNodeOutputs_52; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_107 = io_selectInput_88 ? io_dataInput_88 : io_dataInput_89; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_108 = io_selectInput_90 ? io_dataInput_90 : io_dataInput_91; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_53 = selectNodeOutputs_107 ? dataNodeOutputs_107 : dataNodeOutputs_108; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_109 = io_selectInput_92 ? io_dataInput_92 : io_dataInput_93; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_110 = io_selectInput_94 ? io_dataInput_94 : io_dataInput_95; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_54 = selectNodeOutputs_109 ? dataNodeOutputs_109 : dataNodeOutputs_110; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_26 = selectNodeOutputs_53 ? dataNodeOutputs_53 : dataNodeOutputs_54; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_12 = selectNodeOutputs_25 ? dataNodeOutputs_25 : dataNodeOutputs_26; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_5 = selectNodeOutputs_11 ? dataNodeOutputs_11 : dataNodeOutputs_12; // @[GameUtilities.scala 91:34]
  wire  selectNodeOutputs_111 = io_selectInput_96 | io_selectInput_97; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_112 = io_selectInput_98 | io_selectInput_99; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_55 = selectNodeOutputs_111 | selectNodeOutputs_112; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_113 = io_selectInput_100 | io_selectInput_101; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_114 = io_selectInput_102 | io_selectInput_103; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_56 = selectNodeOutputs_113 | selectNodeOutputs_114; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_27 = selectNodeOutputs_55 | selectNodeOutputs_56; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_115 = io_selectInput_104 | io_selectInput_105; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_116 = io_selectInput_106 | io_selectInput_107; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_57 = selectNodeOutputs_115 | selectNodeOutputs_116; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_117 = io_selectInput_108 | io_selectInput_109; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_118 = io_selectInput_110 | io_selectInput_111; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_58 = selectNodeOutputs_117 | selectNodeOutputs_118; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_28 = selectNodeOutputs_57 | selectNodeOutputs_58; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_13 = selectNodeOutputs_27 | selectNodeOutputs_28; // @[GameUtilities.scala 92:54]
  wire [6:0] dataNodeOutputs_111 = io_selectInput_96 ? io_dataInput_96 : io_dataInput_97; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_112 = io_selectInput_98 ? io_dataInput_98 : io_dataInput_99; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_55 = selectNodeOutputs_111 ? dataNodeOutputs_111 : dataNodeOutputs_112; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_113 = io_selectInput_100 ? io_dataInput_100 : io_dataInput_101; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_114 = io_selectInput_102 ? io_dataInput_102 : io_dataInput_103; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_56 = selectNodeOutputs_113 ? dataNodeOutputs_113 : dataNodeOutputs_114; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_27 = selectNodeOutputs_55 ? dataNodeOutputs_55 : dataNodeOutputs_56; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_115 = io_selectInput_104 ? io_dataInput_104 : io_dataInput_105; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_116 = io_selectInput_106 ? io_dataInput_106 : io_dataInput_107; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_57 = selectNodeOutputs_115 ? dataNodeOutputs_115 : dataNodeOutputs_116; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_117 = io_selectInput_108 ? io_dataInput_108 : io_dataInput_109; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_118 = io_selectInput_110 ? io_dataInput_110 : io_dataInput_111; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_58 = selectNodeOutputs_117 ? dataNodeOutputs_117 : dataNodeOutputs_118; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_28 = selectNodeOutputs_57 ? dataNodeOutputs_57 : dataNodeOutputs_58; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_13 = selectNodeOutputs_27 ? dataNodeOutputs_27 : dataNodeOutputs_28; // @[GameUtilities.scala 91:34]
  wire  selectNodeOutputs_119 = io_selectInput_112 | io_selectInput_113; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_120 = io_selectInput_114 | io_selectInput_115; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_59 = selectNodeOutputs_119 | selectNodeOutputs_120; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_121 = io_selectInput_116 | io_selectInput_117; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_122 = io_selectInput_118 | io_selectInput_119; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_60 = selectNodeOutputs_121 | selectNodeOutputs_122; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_29 = selectNodeOutputs_59 | selectNodeOutputs_60; // @[GameUtilities.scala 92:54]
  wire [6:0] dataNodeOutputs_119 = io_selectInput_112 ? io_dataInput_112 : io_dataInput_113; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_120 = io_selectInput_114 ? io_dataInput_114 : io_dataInput_115; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_59 = selectNodeOutputs_119 ? dataNodeOutputs_119 : dataNodeOutputs_120; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_121 = io_selectInput_116 ? io_dataInput_116 : io_dataInput_117; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_122 = io_selectInput_118 ? io_dataInput_118 : io_dataInput_119; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_60 = selectNodeOutputs_121 ? dataNodeOutputs_121 : dataNodeOutputs_122; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_29 = selectNodeOutputs_59 ? dataNodeOutputs_59 : dataNodeOutputs_60; // @[GameUtilities.scala 91:34]
  wire  selectNodeOutputs_123 = io_selectInput_120 | io_selectInput_121; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_124 = io_selectInput_122 | io_selectInput_123; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_61 = selectNodeOutputs_123 | selectNodeOutputs_124; // @[GameUtilities.scala 92:54]
  wire [6:0] dataNodeOutputs_123 = io_selectInput_120 ? io_dataInput_120 : io_dataInput_121; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_124 = io_selectInput_122 ? io_dataInput_122 : io_dataInput_123; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_61 = selectNodeOutputs_123 ? dataNodeOutputs_123 : dataNodeOutputs_124; // @[GameUtilities.scala 91:34]
  wire  selectNodeOutputs_125 = io_selectInput_124 | io_selectInput_125; // @[GameUtilities.scala 92:54]
  wire [6:0] dataNodeOutputs_125 = io_selectInput_124 ? io_dataInput_124 : io_dataInput_125; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_126 = io_selectInput_126 ? io_dataInput_126 : io_dataInput_127; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_62 = selectNodeOutputs_125 ? dataNodeOutputs_125 : dataNodeOutputs_126; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_30 = selectNodeOutputs_61 ? dataNodeOutputs_61 : dataNodeOutputs_62; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_14 = selectNodeOutputs_29 ? dataNodeOutputs_29 : dataNodeOutputs_30; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_6 = selectNodeOutputs_13 ? dataNodeOutputs_13 : dataNodeOutputs_14; // @[GameUtilities.scala 91:34]
  wire [6:0] dataNodeOutputs_2 = selectNodeOutputs_5 ? dataNodeOutputs_5 : dataNodeOutputs_6; // @[GameUtilities.scala 91:34]
  wire  selectNodeOutputs_126 = io_selectInput_126 | io_selectInput_127; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_62 = selectNodeOutputs_125 | selectNodeOutputs_126; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_30 = selectNodeOutputs_61 | selectNodeOutputs_62; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_14 = selectNodeOutputs_29 | selectNodeOutputs_30; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_6 = selectNodeOutputs_13 | selectNodeOutputs_14; // @[GameUtilities.scala 92:54]
  wire  selectNodeOutputs_2 = selectNodeOutputs_5 | selectNodeOutputs_6; // @[GameUtilities.scala 92:54]
  wire [6:0] indexNodeOutputs_63 = io_selectInput_0 ? 7'h0 : 7'h1; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_64 = io_selectInput_2 ? 7'h2 : 7'h3; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_31 = selectNodeOutputs_63 ? indexNodeOutputs_63 : indexNodeOutputs_64; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_65 = io_selectInput_4 ? 7'h4 : 7'h5; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_66 = io_selectInput_6 ? 7'h6 : 7'h7; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_32 = selectNodeOutputs_65 ? indexNodeOutputs_65 : indexNodeOutputs_66; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_15 = selectNodeOutputs_31 ? indexNodeOutputs_31 : indexNodeOutputs_32; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_67 = io_selectInput_8 ? 7'h8 : 7'h9; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_68 = io_selectInput_10 ? 7'ha : 7'hb; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_33 = selectNodeOutputs_67 ? indexNodeOutputs_67 : indexNodeOutputs_68; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_69 = io_selectInput_12 ? 7'hc : 7'hd; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_70 = io_selectInput_14 ? 7'he : 7'hf; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_34 = selectNodeOutputs_69 ? indexNodeOutputs_69 : indexNodeOutputs_70; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_16 = selectNodeOutputs_33 ? indexNodeOutputs_33 : indexNodeOutputs_34; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_7 = selectNodeOutputs_15 ? indexNodeOutputs_15 : indexNodeOutputs_16; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_71 = io_selectInput_16 ? 7'h10 : 7'h11; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_72 = io_selectInput_18 ? 7'h12 : 7'h13; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_35 = selectNodeOutputs_71 ? indexNodeOutputs_71 : indexNodeOutputs_72; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_73 = io_selectInput_20 ? 7'h14 : 7'h15; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_74 = io_selectInput_22 ? 7'h16 : 7'h17; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_36 = selectNodeOutputs_73 ? indexNodeOutputs_73 : indexNodeOutputs_74; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_17 = selectNodeOutputs_35 ? indexNodeOutputs_35 : indexNodeOutputs_36; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_75 = io_selectInput_24 ? 7'h18 : 7'h19; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_76 = io_selectInput_26 ? 7'h1a : 7'h1b; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_37 = selectNodeOutputs_75 ? indexNodeOutputs_75 : indexNodeOutputs_76; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_77 = io_selectInput_28 ? 7'h1c : 7'h1d; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_78 = io_selectInput_30 ? 7'h1e : 7'h1f; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_38 = selectNodeOutputs_77 ? indexNodeOutputs_77 : indexNodeOutputs_78; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_18 = selectNodeOutputs_37 ? indexNodeOutputs_37 : indexNodeOutputs_38; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_8 = selectNodeOutputs_17 ? indexNodeOutputs_17 : indexNodeOutputs_18; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_3 = selectNodeOutputs_7 ? indexNodeOutputs_7 : indexNodeOutputs_8; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_79 = io_selectInput_32 ? 7'h20 : 7'h21; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_80 = io_selectInput_34 ? 7'h22 : 7'h23; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_39 = selectNodeOutputs_79 ? indexNodeOutputs_79 : indexNodeOutputs_80; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_81 = io_selectInput_36 ? 7'h24 : 7'h25; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_82 = io_selectInput_38 ? 7'h26 : 7'h27; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_40 = selectNodeOutputs_81 ? indexNodeOutputs_81 : indexNodeOutputs_82; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_19 = selectNodeOutputs_39 ? indexNodeOutputs_39 : indexNodeOutputs_40; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_83 = io_selectInput_40 ? 7'h28 : 7'h29; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_84 = io_selectInput_42 ? 7'h2a : 7'h2b; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_41 = selectNodeOutputs_83 ? indexNodeOutputs_83 : indexNodeOutputs_84; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_85 = io_selectInput_44 ? 7'h2c : 7'h2d; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_86 = io_selectInput_46 ? 7'h2e : 7'h2f; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_42 = selectNodeOutputs_85 ? indexNodeOutputs_85 : indexNodeOutputs_86; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_20 = selectNodeOutputs_41 ? indexNodeOutputs_41 : indexNodeOutputs_42; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_9 = selectNodeOutputs_19 ? indexNodeOutputs_19 : indexNodeOutputs_20; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_87 = io_selectInput_48 ? 7'h30 : 7'h31; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_88 = io_selectInput_50 ? 7'h32 : 7'h33; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_43 = selectNodeOutputs_87 ? indexNodeOutputs_87 : indexNodeOutputs_88; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_89 = io_selectInput_52 ? 7'h34 : 7'h35; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_90 = io_selectInput_54 ? 7'h36 : 7'h37; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_44 = selectNodeOutputs_89 ? indexNodeOutputs_89 : indexNodeOutputs_90; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_21 = selectNodeOutputs_43 ? indexNodeOutputs_43 : indexNodeOutputs_44; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_91 = io_selectInput_56 ? 7'h38 : 7'h39; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_92 = io_selectInput_58 ? 7'h3a : 7'h3b; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_45 = selectNodeOutputs_91 ? indexNodeOutputs_91 : indexNodeOutputs_92; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_93 = io_selectInput_60 ? 7'h3c : 7'h3d; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_94 = io_selectInput_62 ? 7'h3e : 7'h3f; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_46 = selectNodeOutputs_93 ? indexNodeOutputs_93 : indexNodeOutputs_94; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_22 = selectNodeOutputs_45 ? indexNodeOutputs_45 : indexNodeOutputs_46; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_10 = selectNodeOutputs_21 ? indexNodeOutputs_21 : indexNodeOutputs_22; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_4 = selectNodeOutputs_9 ? indexNodeOutputs_9 : indexNodeOutputs_10; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_1 = selectNodeOutputs_3 ? indexNodeOutputs_3 : indexNodeOutputs_4; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_95 = io_selectInput_64 ? 7'h40 : 7'h41; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_96 = io_selectInput_66 ? 7'h42 : 7'h43; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_47 = selectNodeOutputs_95 ? indexNodeOutputs_95 : indexNodeOutputs_96; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_97 = io_selectInput_68 ? 7'h44 : 7'h45; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_98 = io_selectInput_70 ? 7'h46 : 7'h47; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_48 = selectNodeOutputs_97 ? indexNodeOutputs_97 : indexNodeOutputs_98; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_23 = selectNodeOutputs_47 ? indexNodeOutputs_47 : indexNodeOutputs_48; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_99 = io_selectInput_72 ? 7'h48 : 7'h49; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_100 = io_selectInput_74 ? 7'h4a : 7'h4b; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_49 = selectNodeOutputs_99 ? indexNodeOutputs_99 : indexNodeOutputs_100; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_101 = io_selectInput_76 ? 7'h4c : 7'h4d; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_102 = io_selectInput_78 ? 7'h4e : 7'h4f; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_50 = selectNodeOutputs_101 ? indexNodeOutputs_101 : indexNodeOutputs_102; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_24 = selectNodeOutputs_49 ? indexNodeOutputs_49 : indexNodeOutputs_50; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_11 = selectNodeOutputs_23 ? indexNodeOutputs_23 : indexNodeOutputs_24; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_103 = io_selectInput_80 ? 7'h50 : 7'h51; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_104 = io_selectInput_82 ? 7'h52 : 7'h53; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_51 = selectNodeOutputs_103 ? indexNodeOutputs_103 : indexNodeOutputs_104; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_105 = io_selectInput_84 ? 7'h54 : 7'h55; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_106 = io_selectInput_86 ? 7'h56 : 7'h57; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_52 = selectNodeOutputs_105 ? indexNodeOutputs_105 : indexNodeOutputs_106; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_25 = selectNodeOutputs_51 ? indexNodeOutputs_51 : indexNodeOutputs_52; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_107 = io_selectInput_88 ? 7'h58 : 7'h59; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_108 = io_selectInput_90 ? 7'h5a : 7'h5b; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_53 = selectNodeOutputs_107 ? indexNodeOutputs_107 : indexNodeOutputs_108; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_109 = io_selectInput_92 ? 7'h5c : 7'h5d; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_110 = io_selectInput_94 ? 7'h5e : 7'h5f; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_54 = selectNodeOutputs_109 ? indexNodeOutputs_109 : indexNodeOutputs_110; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_26 = selectNodeOutputs_53 ? indexNodeOutputs_53 : indexNodeOutputs_54; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_12 = selectNodeOutputs_25 ? indexNodeOutputs_25 : indexNodeOutputs_26; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_5 = selectNodeOutputs_11 ? indexNodeOutputs_11 : indexNodeOutputs_12; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_111 = io_selectInput_96 ? 7'h60 : 7'h61; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_112 = io_selectInput_98 ? 7'h62 : 7'h63; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_55 = selectNodeOutputs_111 ? indexNodeOutputs_111 : indexNodeOutputs_112; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_113 = io_selectInput_100 ? 7'h64 : 7'h65; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_114 = io_selectInput_102 ? 7'h66 : 7'h67; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_56 = selectNodeOutputs_113 ? indexNodeOutputs_113 : indexNodeOutputs_114; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_27 = selectNodeOutputs_55 ? indexNodeOutputs_55 : indexNodeOutputs_56; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_115 = io_selectInput_104 ? 7'h68 : 7'h69; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_116 = io_selectInput_106 ? 7'h6a : 7'h6b; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_57 = selectNodeOutputs_115 ? indexNodeOutputs_115 : indexNodeOutputs_116; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_117 = io_selectInput_108 ? 7'h6c : 7'h6d; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_118 = io_selectInput_110 ? 7'h6e : 7'h6f; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_58 = selectNodeOutputs_117 ? indexNodeOutputs_117 : indexNodeOutputs_118; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_28 = selectNodeOutputs_57 ? indexNodeOutputs_57 : indexNodeOutputs_58; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_13 = selectNodeOutputs_27 ? indexNodeOutputs_27 : indexNodeOutputs_28; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_119 = io_selectInput_112 ? 7'h70 : 7'h71; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_120 = io_selectInput_114 ? 7'h72 : 7'h73; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_59 = selectNodeOutputs_119 ? indexNodeOutputs_119 : indexNodeOutputs_120; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_121 = io_selectInput_116 ? 7'h74 : 7'h75; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_122 = io_selectInput_118 ? 7'h76 : 7'h77; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_60 = selectNodeOutputs_121 ? indexNodeOutputs_121 : indexNodeOutputs_122; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_29 = selectNodeOutputs_59 ? indexNodeOutputs_59 : indexNodeOutputs_60; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_123 = io_selectInput_120 ? 7'h78 : 7'h79; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_124 = io_selectInput_122 ? 7'h7a : 7'h7b; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_61 = selectNodeOutputs_123 ? indexNodeOutputs_123 : indexNodeOutputs_124; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_125 = io_selectInput_124 ? 7'h7c : 7'h7d; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_126 = io_selectInput_126 ? 7'h7e : 7'h7f; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_62 = selectNodeOutputs_125 ? indexNodeOutputs_125 : indexNodeOutputs_126; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_30 = selectNodeOutputs_61 ? indexNodeOutputs_61 : indexNodeOutputs_62; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_14 = selectNodeOutputs_29 ? indexNodeOutputs_29 : indexNodeOutputs_30; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_6 = selectNodeOutputs_13 ? indexNodeOutputs_13 : indexNodeOutputs_14; // @[GameUtilities.scala 93:35]
  wire [6:0] indexNodeOutputs_2 = selectNodeOutputs_5 ? indexNodeOutputs_5 : indexNodeOutputs_6; // @[GameUtilities.scala 93:35]
  assign io_dataOutput = selectNodeOutputs_1 ? dataNodeOutputs_1 : dataNodeOutputs_2; // @[GameUtilities.scala 77:17]
  assign io_selectOutput = selectNodeOutputs_1 | selectNodeOutputs_2; // @[GameUtilities.scala 78:19]
  assign io_indexOutput = selectNodeOutputs_1 ? indexNodeOutputs_1 : indexNodeOutputs_2; // @[GameUtilities.scala 79:18]
endmodule
module SpriteBlender(
  input        clock,
  input  [5:0] io_pixelColorBack,
  input        io_spriteVisibleReg_0,
  input        io_spriteVisibleReg_1,
  input        io_spriteVisibleReg_2,
  input        io_spriteVisibleReg_3,
  input        io_spriteVisibleReg_4,
  input        io_spriteVisibleReg_5,
  input        io_spriteVisibleReg_6,
  input        io_spriteVisibleReg_7,
  input        io_spriteVisibleReg_8,
  input        io_spriteVisibleReg_9,
  input        io_spriteVisibleReg_10,
  input        io_spriteVisibleReg_11,
  input        io_spriteVisibleReg_12,
  input        io_spriteVisibleReg_13,
  input        io_spriteVisibleReg_14,
  input        io_spriteVisibleReg_15,
  input        io_spriteVisibleReg_16,
  input        io_spriteVisibleReg_17,
  input        io_spriteVisibleReg_18,
  input        io_spriteVisibleReg_19,
  input        io_spriteVisibleReg_20,
  input        io_spriteVisibleReg_21,
  input        io_spriteVisibleReg_22,
  input        io_spriteVisibleReg_23,
  input        io_spriteVisibleReg_24,
  input        io_spriteVisibleReg_25,
  input        io_spriteVisibleReg_26,
  input        io_spriteVisibleReg_27,
  input        io_spriteVisibleReg_28,
  input        io_spriteVisibleReg_29,
  input        io_spriteVisibleReg_30,
  input        io_spriteVisibleReg_31,
  input        io_spriteVisibleReg_32,
  input        io_spriteVisibleReg_33,
  input        io_spriteVisibleReg_41,
  input        io_spriteVisibleReg_42,
  input        io_spriteVisibleReg_43,
  input        io_spriteVisibleReg_44,
  input        io_spriteVisibleReg_45,
  input        io_spriteVisibleReg_46,
  input        io_spriteVisibleReg_47,
  input        io_spriteVisibleReg_48,
  input        io_spriteVisibleReg_49,
  input        io_spriteVisibleReg_50,
  input        io_spriteVisibleReg_51,
  input        io_spriteVisibleReg_55,
  input        io_spriteVisibleReg_56,
  input        io_spriteVisibleReg_57,
  input        io_spriteVisibleReg_61,
  input        io_spriteVisibleReg_62,
  input        io_spriteVisibleReg_63,
  input        io_spriteVisibleReg_64,
  input        io_spriteVisibleReg_65,
  input        io_spriteVisibleReg_66,
  input        io_spriteVisibleReg_70,
  input        io_spriteVisibleReg_71,
  input        io_spriteVisibleReg_72,
  input        io_inSprite_0,
  input        io_inSprite_1,
  input        io_inSprite_2,
  input        io_inSprite_3,
  input        io_inSprite_4,
  input        io_inSprite_5,
  input        io_inSprite_6,
  input        io_inSprite_7,
  input        io_inSprite_8,
  input        io_inSprite_9,
  input        io_inSprite_10,
  input        io_inSprite_11,
  input        io_inSprite_12,
  input        io_inSprite_13,
  input        io_inSprite_14,
  input        io_inSprite_15,
  input        io_inSprite_16,
  input        io_inSprite_17,
  input        io_inSprite_18,
  input        io_inSprite_19,
  input        io_inSprite_20,
  input        io_inSprite_21,
  input        io_inSprite_22,
  input        io_inSprite_23,
  input        io_inSprite_24,
  input        io_inSprite_25,
  input        io_inSprite_26,
  input        io_inSprite_27,
  input        io_inSprite_28,
  input        io_inSprite_29,
  input        io_inSprite_30,
  input        io_inSprite_31,
  input        io_inSprite_32,
  input        io_inSprite_33,
  input        io_inSprite_34,
  input        io_inSprite_35,
  input        io_inSprite_36,
  input        io_inSprite_37,
  input        io_inSprite_38,
  input        io_inSprite_39,
  input        io_inSprite_40,
  input        io_inSprite_41,
  input        io_inSprite_42,
  input        io_inSprite_43,
  input        io_inSprite_44,
  input        io_inSprite_45,
  input        io_inSprite_46,
  input        io_inSprite_47,
  input        io_inSprite_48,
  input        io_inSprite_49,
  input        io_inSprite_50,
  input        io_inSprite_51,
  input        io_inSprite_52,
  input        io_inSprite_53,
  input        io_inSprite_54,
  input        io_inSprite_55,
  input        io_inSprite_56,
  input        io_inSprite_57,
  input        io_inSprite_58,
  input        io_inSprite_59,
  input        io_inSprite_60,
  input        io_inSprite_61,
  input        io_inSprite_62,
  input        io_inSprite_63,
  input        io_inSprite_64,
  input        io_inSprite_65,
  input        io_inSprite_66,
  input        io_inSprite_67,
  input        io_inSprite_68,
  input        io_inSprite_69,
  input        io_inSprite_70,
  input        io_inSprite_71,
  input        io_inSprite_72,
  input        io_inSprite_73,
  input        io_inSprite_74,
  input        io_inSprite_75,
  input        io_inSprite_76,
  input        io_inSprite_77,
  input        io_inSprite_78,
  input        io_inSprite_79,
  input        io_inSprite_80,
  input        io_inSprite_81,
  input        io_inSprite_82,
  input        io_inSprite_83,
  input        io_inSprite_84,
  input        io_inSprite_85,
  input        io_inSprite_86,
  input        io_inSprite_87,
  input        io_inSprite_88,
  input        io_inSprite_89,
  input        io_inSprite_90,
  input        io_inSprite_91,
  input        io_inSprite_92,
  input        io_inSprite_93,
  input        io_inSprite_94,
  input        io_inSprite_95,
  input        io_inSprite_96,
  input        io_inSprite_97,
  input        io_inSprite_98,
  input        io_inSprite_99,
  input        io_inSprite_100,
  input        io_inSprite_101,
  input        io_inSprite_102,
  input        io_inSprite_103,
  input        io_inSprite_104,
  input        io_inSprite_105,
  input        io_inSprite_106,
  input        io_inSprite_107,
  input        io_inSprite_108,
  input        io_inSprite_109,
  input        io_inSprite_110,
  input        io_inSprite_111,
  input        io_inSprite_112,
  input        io_inSprite_113,
  input        io_inSprite_114,
  input        io_inSprite_115,
  input        io_inSprite_116,
  input        io_inSprite_117,
  input        io_inSprite_118,
  input        io_inSprite_119,
  input        io_inSprite_120,
  input        io_inSprite_121,
  input        io_inSprite_122,
  input        io_inSprite_123,
  input        io_inSprite_124,
  input        io_inSprite_125,
  input        io_inSprite_126,
  input        io_inSprite_127,
  input  [6:0] io_datareader_0,
  input  [6:0] io_datareader_1,
  input  [6:0] io_datareader_2,
  input  [6:0] io_datareader_3,
  input  [6:0] io_datareader_4,
  input  [6:0] io_datareader_5,
  input  [6:0] io_datareader_6,
  input  [6:0] io_datareader_7,
  input  [6:0] io_datareader_8,
  input  [6:0] io_datareader_9,
  input  [6:0] io_datareader_10,
  input  [6:0] io_datareader_11,
  input  [6:0] io_datareader_12,
  input  [6:0] io_datareader_13,
  input  [6:0] io_datareader_14,
  input  [6:0] io_datareader_15,
  input  [6:0] io_datareader_16,
  input  [6:0] io_datareader_17,
  input  [6:0] io_datareader_18,
  input  [6:0] io_datareader_19,
  input  [6:0] io_datareader_20,
  input  [6:0] io_datareader_21,
  input  [6:0] io_datareader_22,
  input  [6:0] io_datareader_23,
  input  [6:0] io_datareader_24,
  input  [6:0] io_datareader_25,
  input  [6:0] io_datareader_26,
  input  [6:0] io_datareader_27,
  input  [6:0] io_datareader_28,
  input  [6:0] io_datareader_29,
  input  [6:0] io_datareader_30,
  input  [6:0] io_datareader_31,
  input  [6:0] io_datareader_32,
  input  [6:0] io_datareader_33,
  input  [6:0] io_datareader_34,
  input  [6:0] io_datareader_35,
  input  [6:0] io_datareader_36,
  input  [6:0] io_datareader_37,
  input  [6:0] io_datareader_38,
  input  [6:0] io_datareader_39,
  input  [6:0] io_datareader_40,
  input  [6:0] io_datareader_41,
  input  [6:0] io_datareader_42,
  input  [6:0] io_datareader_43,
  input  [6:0] io_datareader_44,
  input  [6:0] io_datareader_45,
  input  [6:0] io_datareader_46,
  input  [6:0] io_datareader_47,
  input  [6:0] io_datareader_48,
  input  [6:0] io_datareader_49,
  input  [6:0] io_datareader_50,
  input  [6:0] io_datareader_51,
  input  [6:0] io_datareader_52,
  input  [6:0] io_datareader_53,
  input  [6:0] io_datareader_54,
  input  [6:0] io_datareader_55,
  input  [6:0] io_datareader_56,
  input  [6:0] io_datareader_57,
  input  [6:0] io_datareader_58,
  input  [6:0] io_datareader_59,
  input  [6:0] io_datareader_60,
  input  [6:0] io_datareader_61,
  input  [6:0] io_datareader_62,
  input  [6:0] io_datareader_63,
  input  [6:0] io_datareader_64,
  input  [6:0] io_datareader_65,
  input  [6:0] io_datareader_66,
  input  [6:0] io_datareader_67,
  input  [6:0] io_datareader_68,
  input  [6:0] io_datareader_69,
  input  [6:0] io_datareader_70,
  input  [6:0] io_datareader_71,
  input  [6:0] io_datareader_72,
  input  [6:0] io_datareader_73,
  input  [6:0] io_datareader_74,
  input  [6:0] io_datareader_75,
  input  [6:0] io_datareader_76,
  input  [6:0] io_datareader_77,
  input  [6:0] io_datareader_78,
  input  [6:0] io_datareader_79,
  input  [6:0] io_datareader_80,
  input  [6:0] io_datareader_81,
  input  [6:0] io_datareader_82,
  input  [6:0] io_datareader_83,
  input  [6:0] io_datareader_84,
  input  [6:0] io_datareader_85,
  input  [6:0] io_datareader_86,
  input  [6:0] io_datareader_87,
  input  [6:0] io_datareader_88,
  input  [6:0] io_datareader_89,
  input  [6:0] io_datareader_90,
  input  [6:0] io_datareader_91,
  input  [6:0] io_datareader_92,
  input  [6:0] io_datareader_93,
  input  [6:0] io_datareader_94,
  input  [6:0] io_datareader_95,
  input  [6:0] io_datareader_96,
  input  [6:0] io_datareader_97,
  input  [6:0] io_datareader_98,
  input  [6:0] io_datareader_99,
  input  [6:0] io_datareader_100,
  input  [6:0] io_datareader_101,
  input  [6:0] io_datareader_102,
  input  [6:0] io_datareader_103,
  input  [6:0] io_datareader_104,
  input  [6:0] io_datareader_105,
  input  [6:0] io_datareader_106,
  input  [6:0] io_datareader_107,
  input  [6:0] io_datareader_108,
  input  [6:0] io_datareader_109,
  input  [6:0] io_datareader_110,
  input  [6:0] io_datareader_111,
  input  [6:0] io_datareader_112,
  input  [6:0] io_datareader_113,
  input  [6:0] io_datareader_114,
  input  [6:0] io_datareader_115,
  input  [6:0] io_datareader_116,
  input  [6:0] io_datareader_117,
  input  [6:0] io_datareader_118,
  input  [6:0] io_datareader_119,
  input  [6:0] io_datareader_120,
  input  [6:0] io_datareader_121,
  input  [6:0] io_datareader_122,
  input  [6:0] io_datareader_123,
  input  [6:0] io_datareader_124,
  input  [6:0] io_datareader_125,
  input  [6:0] io_datareader_126,
  input  [6:0] io_datareader_127,
  output [3:0] io_vgaRed,
  output [3:0] io_vgaGreen,
  output [3:0] io_vgaBlue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_0; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_1; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_2; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_3; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_4; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_5; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_6; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_7; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_8; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_9; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_10; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_11; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_12; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_13; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_14; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_15; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_16; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_17; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_18; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_19; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_20; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_21; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_22; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_23; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_24; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_25; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_26; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_27; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_28; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_29; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_30; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_31; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_32; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_33; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_34; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_35; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_36; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_37; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_38; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_39; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_40; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_41; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_42; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_43; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_44; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_45; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_46; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_47; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_48; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_49; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_50; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_51; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_52; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_53; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_54; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_55; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_56; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_57; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_58; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_59; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_60; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_61; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_62; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_63; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_64; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_65; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_66; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_67; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_68; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_69; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_70; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_71; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_72; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_73; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_74; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_75; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_76; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_77; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_78; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_79; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_80; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_81; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_82; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_83; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_84; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_85; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_86; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_87; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_88; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_89; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_90; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_91; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_92; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_93; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_94; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_95; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_96; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_97; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_98; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_99; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_100; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_101; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_102; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_103; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_104; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_105; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_106; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_107; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_108; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_109; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_110; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_111; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_112; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_113; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_114; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_115; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_116; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_117; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_118; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_119; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_120; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_121; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_122; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_123; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_124; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_125; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_126; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataInput_127; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_0; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_1; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_2; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_3; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_4; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_5; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_6; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_7; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_8; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_9; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_10; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_11; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_12; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_13; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_14; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_15; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_16; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_17; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_18; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_19; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_20; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_21; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_22; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_23; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_24; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_25; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_26; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_27; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_28; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_29; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_30; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_31; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_32; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_33; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_34; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_35; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_36; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_37; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_38; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_39; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_40; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_41; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_42; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_43; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_44; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_45; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_46; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_47; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_48; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_49; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_50; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_51; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_52; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_53; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_54; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_55; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_56; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_57; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_58; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_59; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_60; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_61; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_62; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_63; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_64; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_65; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_66; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_67; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_68; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_69; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_70; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_71; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_72; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_73; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_74; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_75; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_76; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_77; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_78; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_79; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_80; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_81; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_82; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_83; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_84; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_85; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_86; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_87; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_88; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_89; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_90; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_91; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_92; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_93; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_94; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_95; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_96; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_97; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_98; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_99; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_100; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_101; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_102; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_103; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_104; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_105; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_106; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_107; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_108; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_109; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_110; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_111; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_112; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_113; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_114; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_115; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_116; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_117; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_118; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_119; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_120; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_121; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_122; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_123; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_124; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_125; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_126; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectInput_127; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_dataOutput; // @[SpriteBlender.scala 33:44]
  wire  multiHotPriortyReductionTree_io_selectOutput; // @[SpriteBlender.scala 33:44]
  wire [6:0] multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 33:44]
  reg [5:0] _T; // @[SpriteBlender.scala 23:42]
  reg [5:0] pixelColorBackReg; // @[SpriteBlender.scala 23:34]
  reg  _T_3_0; // @[GameUtilities.scala 21:24]
  reg  _T_3_1; // @[GameUtilities.scala 21:24]
  reg  _T_4_0; // @[GameUtilities.scala 21:24]
  reg  _T_4_1; // @[GameUtilities.scala 21:24]
  wire  _T_5 = _T_3_0 & _T_4_0; // @[SpriteBlender.scala 40:43]
  wire  _T_7 = ~io_datareader_0[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_11_0; // @[GameUtilities.scala 21:24]
  reg  _T_11_1; // @[GameUtilities.scala 21:24]
  reg  _T_12_0; // @[GameUtilities.scala 21:24]
  reg  _T_12_1; // @[GameUtilities.scala 21:24]
  wire  _T_13 = _T_11_0 & _T_12_0; // @[SpriteBlender.scala 40:43]
  wire  _T_15 = ~io_datareader_1[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_19_0; // @[GameUtilities.scala 21:24]
  reg  _T_19_1; // @[GameUtilities.scala 21:24]
  reg  _T_20_0; // @[GameUtilities.scala 21:24]
  reg  _T_20_1; // @[GameUtilities.scala 21:24]
  wire  _T_21 = _T_19_0 & _T_20_0; // @[SpriteBlender.scala 40:43]
  wire  _T_23 = ~io_datareader_2[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_27_0; // @[GameUtilities.scala 21:24]
  reg  _T_27_1; // @[GameUtilities.scala 21:24]
  reg  _T_28_0; // @[GameUtilities.scala 21:24]
  reg  _T_28_1; // @[GameUtilities.scala 21:24]
  wire  _T_29 = _T_27_0 & _T_28_0; // @[SpriteBlender.scala 40:43]
  wire  _T_31 = ~io_datareader_3[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_35_0; // @[GameUtilities.scala 21:24]
  reg  _T_35_1; // @[GameUtilities.scala 21:24]
  reg  _T_36_0; // @[GameUtilities.scala 21:24]
  reg  _T_36_1; // @[GameUtilities.scala 21:24]
  wire  _T_37 = _T_35_0 & _T_36_0; // @[SpriteBlender.scala 40:43]
  wire  _T_39 = ~io_datareader_4[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_43_0; // @[GameUtilities.scala 21:24]
  reg  _T_43_1; // @[GameUtilities.scala 21:24]
  reg  _T_44_0; // @[GameUtilities.scala 21:24]
  reg  _T_44_1; // @[GameUtilities.scala 21:24]
  wire  _T_45 = _T_43_0 & _T_44_0; // @[SpriteBlender.scala 40:43]
  wire  _T_47 = ~io_datareader_5[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_51_0; // @[GameUtilities.scala 21:24]
  reg  _T_51_1; // @[GameUtilities.scala 21:24]
  reg  _T_52_0; // @[GameUtilities.scala 21:24]
  reg  _T_52_1; // @[GameUtilities.scala 21:24]
  wire  _T_53 = _T_51_0 & _T_52_0; // @[SpriteBlender.scala 40:43]
  wire  _T_55 = ~io_datareader_6[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_59_0; // @[GameUtilities.scala 21:24]
  reg  _T_59_1; // @[GameUtilities.scala 21:24]
  reg  _T_60_0; // @[GameUtilities.scala 21:24]
  reg  _T_60_1; // @[GameUtilities.scala 21:24]
  wire  _T_61 = _T_59_0 & _T_60_0; // @[SpriteBlender.scala 40:43]
  wire  _T_63 = ~io_datareader_7[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_67_0; // @[GameUtilities.scala 21:24]
  reg  _T_67_1; // @[GameUtilities.scala 21:24]
  reg  _T_68_0; // @[GameUtilities.scala 21:24]
  reg  _T_68_1; // @[GameUtilities.scala 21:24]
  wire  _T_69 = _T_67_0 & _T_68_0; // @[SpriteBlender.scala 40:43]
  wire  _T_71 = ~io_datareader_8[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_75_0; // @[GameUtilities.scala 21:24]
  reg  _T_75_1; // @[GameUtilities.scala 21:24]
  reg  _T_76_0; // @[GameUtilities.scala 21:24]
  reg  _T_76_1; // @[GameUtilities.scala 21:24]
  wire  _T_77 = _T_75_0 & _T_76_0; // @[SpriteBlender.scala 40:43]
  wire  _T_79 = ~io_datareader_9[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_83_0; // @[GameUtilities.scala 21:24]
  reg  _T_83_1; // @[GameUtilities.scala 21:24]
  reg  _T_84_0; // @[GameUtilities.scala 21:24]
  reg  _T_84_1; // @[GameUtilities.scala 21:24]
  wire  _T_85 = _T_83_0 & _T_84_0; // @[SpriteBlender.scala 40:43]
  wire  _T_87 = ~io_datareader_10[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_91_0; // @[GameUtilities.scala 21:24]
  reg  _T_91_1; // @[GameUtilities.scala 21:24]
  reg  _T_92_0; // @[GameUtilities.scala 21:24]
  reg  _T_92_1; // @[GameUtilities.scala 21:24]
  wire  _T_93 = _T_91_0 & _T_92_0; // @[SpriteBlender.scala 40:43]
  wire  _T_95 = ~io_datareader_11[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_99_0; // @[GameUtilities.scala 21:24]
  reg  _T_99_1; // @[GameUtilities.scala 21:24]
  reg  _T_100_0; // @[GameUtilities.scala 21:24]
  reg  _T_100_1; // @[GameUtilities.scala 21:24]
  wire  _T_101 = _T_99_0 & _T_100_0; // @[SpriteBlender.scala 40:43]
  wire  _T_103 = ~io_datareader_12[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_107_0; // @[GameUtilities.scala 21:24]
  reg  _T_107_1; // @[GameUtilities.scala 21:24]
  reg  _T_108_0; // @[GameUtilities.scala 21:24]
  reg  _T_108_1; // @[GameUtilities.scala 21:24]
  wire  _T_109 = _T_107_0 & _T_108_0; // @[SpriteBlender.scala 40:43]
  wire  _T_111 = ~io_datareader_13[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_115_0; // @[GameUtilities.scala 21:24]
  reg  _T_115_1; // @[GameUtilities.scala 21:24]
  reg  _T_116_0; // @[GameUtilities.scala 21:24]
  reg  _T_116_1; // @[GameUtilities.scala 21:24]
  wire  _T_117 = _T_115_0 & _T_116_0; // @[SpriteBlender.scala 40:43]
  wire  _T_119 = ~io_datareader_14[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_123_0; // @[GameUtilities.scala 21:24]
  reg  _T_123_1; // @[GameUtilities.scala 21:24]
  reg  _T_124_0; // @[GameUtilities.scala 21:24]
  reg  _T_124_1; // @[GameUtilities.scala 21:24]
  wire  _T_125 = _T_123_0 & _T_124_0; // @[SpriteBlender.scala 40:43]
  wire  _T_127 = ~io_datareader_15[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_131_0; // @[GameUtilities.scala 21:24]
  reg  _T_131_1; // @[GameUtilities.scala 21:24]
  reg  _T_132_0; // @[GameUtilities.scala 21:24]
  reg  _T_132_1; // @[GameUtilities.scala 21:24]
  wire  _T_133 = _T_131_0 & _T_132_0; // @[SpriteBlender.scala 40:43]
  wire  _T_135 = ~io_datareader_16[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_139_0; // @[GameUtilities.scala 21:24]
  reg  _T_139_1; // @[GameUtilities.scala 21:24]
  reg  _T_140_0; // @[GameUtilities.scala 21:24]
  reg  _T_140_1; // @[GameUtilities.scala 21:24]
  wire  _T_141 = _T_139_0 & _T_140_0; // @[SpriteBlender.scala 40:43]
  wire  _T_143 = ~io_datareader_17[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_147_0; // @[GameUtilities.scala 21:24]
  reg  _T_147_1; // @[GameUtilities.scala 21:24]
  reg  _T_148_0; // @[GameUtilities.scala 21:24]
  reg  _T_148_1; // @[GameUtilities.scala 21:24]
  wire  _T_149 = _T_147_0 & _T_148_0; // @[SpriteBlender.scala 40:43]
  wire  _T_151 = ~io_datareader_18[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_155_0; // @[GameUtilities.scala 21:24]
  reg  _T_155_1; // @[GameUtilities.scala 21:24]
  reg  _T_156_0; // @[GameUtilities.scala 21:24]
  reg  _T_156_1; // @[GameUtilities.scala 21:24]
  wire  _T_157 = _T_155_0 & _T_156_0; // @[SpriteBlender.scala 40:43]
  wire  _T_159 = ~io_datareader_19[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_163_0; // @[GameUtilities.scala 21:24]
  reg  _T_163_1; // @[GameUtilities.scala 21:24]
  reg  _T_164_0; // @[GameUtilities.scala 21:24]
  reg  _T_164_1; // @[GameUtilities.scala 21:24]
  wire  _T_165 = _T_163_0 & _T_164_0; // @[SpriteBlender.scala 40:43]
  wire  _T_167 = ~io_datareader_20[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_171_0; // @[GameUtilities.scala 21:24]
  reg  _T_171_1; // @[GameUtilities.scala 21:24]
  reg  _T_172_0; // @[GameUtilities.scala 21:24]
  reg  _T_172_1; // @[GameUtilities.scala 21:24]
  wire  _T_173 = _T_171_0 & _T_172_0; // @[SpriteBlender.scala 40:43]
  wire  _T_175 = ~io_datareader_21[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_179_0; // @[GameUtilities.scala 21:24]
  reg  _T_179_1; // @[GameUtilities.scala 21:24]
  reg  _T_180_0; // @[GameUtilities.scala 21:24]
  reg  _T_180_1; // @[GameUtilities.scala 21:24]
  wire  _T_181 = _T_179_0 & _T_180_0; // @[SpriteBlender.scala 40:43]
  wire  _T_183 = ~io_datareader_22[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_187_0; // @[GameUtilities.scala 21:24]
  reg  _T_187_1; // @[GameUtilities.scala 21:24]
  reg  _T_188_0; // @[GameUtilities.scala 21:24]
  reg  _T_188_1; // @[GameUtilities.scala 21:24]
  wire  _T_189 = _T_187_0 & _T_188_0; // @[SpriteBlender.scala 40:43]
  wire  _T_191 = ~io_datareader_23[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_195_0; // @[GameUtilities.scala 21:24]
  reg  _T_195_1; // @[GameUtilities.scala 21:24]
  reg  _T_196_0; // @[GameUtilities.scala 21:24]
  reg  _T_196_1; // @[GameUtilities.scala 21:24]
  wire  _T_197 = _T_195_0 & _T_196_0; // @[SpriteBlender.scala 40:43]
  wire  _T_199 = ~io_datareader_24[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_203_0; // @[GameUtilities.scala 21:24]
  reg  _T_203_1; // @[GameUtilities.scala 21:24]
  reg  _T_204_0; // @[GameUtilities.scala 21:24]
  reg  _T_204_1; // @[GameUtilities.scala 21:24]
  wire  _T_205 = _T_203_0 & _T_204_0; // @[SpriteBlender.scala 40:43]
  wire  _T_207 = ~io_datareader_25[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_211_0; // @[GameUtilities.scala 21:24]
  reg  _T_211_1; // @[GameUtilities.scala 21:24]
  reg  _T_212_0; // @[GameUtilities.scala 21:24]
  reg  _T_212_1; // @[GameUtilities.scala 21:24]
  wire  _T_213 = _T_211_0 & _T_212_0; // @[SpriteBlender.scala 40:43]
  wire  _T_215 = ~io_datareader_26[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_219_0; // @[GameUtilities.scala 21:24]
  reg  _T_219_1; // @[GameUtilities.scala 21:24]
  reg  _T_220_0; // @[GameUtilities.scala 21:24]
  reg  _T_220_1; // @[GameUtilities.scala 21:24]
  wire  _T_221 = _T_219_0 & _T_220_0; // @[SpriteBlender.scala 40:43]
  wire  _T_223 = ~io_datareader_27[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_227_0; // @[GameUtilities.scala 21:24]
  reg  _T_227_1; // @[GameUtilities.scala 21:24]
  reg  _T_228_0; // @[GameUtilities.scala 21:24]
  reg  _T_228_1; // @[GameUtilities.scala 21:24]
  wire  _T_229 = _T_227_0 & _T_228_0; // @[SpriteBlender.scala 40:43]
  wire  _T_231 = ~io_datareader_28[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_235_0; // @[GameUtilities.scala 21:24]
  reg  _T_235_1; // @[GameUtilities.scala 21:24]
  reg  _T_236_0; // @[GameUtilities.scala 21:24]
  reg  _T_236_1; // @[GameUtilities.scala 21:24]
  wire  _T_237 = _T_235_0 & _T_236_0; // @[SpriteBlender.scala 40:43]
  wire  _T_239 = ~io_datareader_29[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_243_0; // @[GameUtilities.scala 21:24]
  reg  _T_243_1; // @[GameUtilities.scala 21:24]
  reg  _T_244_0; // @[GameUtilities.scala 21:24]
  reg  _T_244_1; // @[GameUtilities.scala 21:24]
  wire  _T_245 = _T_243_0 & _T_244_0; // @[SpriteBlender.scala 40:43]
  wire  _T_247 = ~io_datareader_30[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_251_0; // @[GameUtilities.scala 21:24]
  reg  _T_251_1; // @[GameUtilities.scala 21:24]
  reg  _T_252_0; // @[GameUtilities.scala 21:24]
  reg  _T_252_1; // @[GameUtilities.scala 21:24]
  wire  _T_253 = _T_251_0 & _T_252_0; // @[SpriteBlender.scala 40:43]
  wire  _T_255 = ~io_datareader_31[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_259_0; // @[GameUtilities.scala 21:24]
  reg  _T_259_1; // @[GameUtilities.scala 21:24]
  reg  _T_260_0; // @[GameUtilities.scala 21:24]
  reg  _T_260_1; // @[GameUtilities.scala 21:24]
  wire  _T_261 = _T_259_0 & _T_260_0; // @[SpriteBlender.scala 40:43]
  wire  _T_263 = ~io_datareader_32[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_267_0; // @[GameUtilities.scala 21:24]
  reg  _T_267_1; // @[GameUtilities.scala 21:24]
  reg  _T_268_0; // @[GameUtilities.scala 21:24]
  reg  _T_268_1; // @[GameUtilities.scala 21:24]
  wire  _T_269 = _T_267_0 & _T_268_0; // @[SpriteBlender.scala 40:43]
  wire  _T_271 = ~io_datareader_33[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_276_0; // @[GameUtilities.scala 21:24]
  reg  _T_276_1; // @[GameUtilities.scala 21:24]
  wire  _T_279 = ~io_datareader_34[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_284_0; // @[GameUtilities.scala 21:24]
  reg  _T_284_1; // @[GameUtilities.scala 21:24]
  wire  _T_287 = ~io_datareader_35[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_292_0; // @[GameUtilities.scala 21:24]
  reg  _T_292_1; // @[GameUtilities.scala 21:24]
  wire  _T_295 = ~io_datareader_36[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_300_0; // @[GameUtilities.scala 21:24]
  reg  _T_300_1; // @[GameUtilities.scala 21:24]
  wire  _T_303 = ~io_datareader_37[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_308_0; // @[GameUtilities.scala 21:24]
  reg  _T_308_1; // @[GameUtilities.scala 21:24]
  wire  _T_311 = ~io_datareader_38[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_316_0; // @[GameUtilities.scala 21:24]
  reg  _T_316_1; // @[GameUtilities.scala 21:24]
  wire  _T_319 = ~io_datareader_39[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_324_0; // @[GameUtilities.scala 21:24]
  reg  _T_324_1; // @[GameUtilities.scala 21:24]
  wire  _T_327 = ~io_datareader_40[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_331_0; // @[GameUtilities.scala 21:24]
  reg  _T_331_1; // @[GameUtilities.scala 21:24]
  reg  _T_332_0; // @[GameUtilities.scala 21:24]
  reg  _T_332_1; // @[GameUtilities.scala 21:24]
  wire  _T_333 = _T_331_0 & _T_332_0; // @[SpriteBlender.scala 40:43]
  wire  _T_335 = ~io_datareader_41[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_339_0; // @[GameUtilities.scala 21:24]
  reg  _T_339_1; // @[GameUtilities.scala 21:24]
  reg  _T_340_0; // @[GameUtilities.scala 21:24]
  reg  _T_340_1; // @[GameUtilities.scala 21:24]
  wire  _T_341 = _T_339_0 & _T_340_0; // @[SpriteBlender.scala 40:43]
  wire  _T_343 = ~io_datareader_42[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_347_0; // @[GameUtilities.scala 21:24]
  reg  _T_347_1; // @[GameUtilities.scala 21:24]
  reg  _T_348_0; // @[GameUtilities.scala 21:24]
  reg  _T_348_1; // @[GameUtilities.scala 21:24]
  wire  _T_349 = _T_347_0 & _T_348_0; // @[SpriteBlender.scala 40:43]
  wire  _T_351 = ~io_datareader_43[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_355_0; // @[GameUtilities.scala 21:24]
  reg  _T_355_1; // @[GameUtilities.scala 21:24]
  reg  _T_356_0; // @[GameUtilities.scala 21:24]
  reg  _T_356_1; // @[GameUtilities.scala 21:24]
  wire  _T_357 = _T_355_0 & _T_356_0; // @[SpriteBlender.scala 40:43]
  wire  _T_359 = ~io_datareader_44[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_363_0; // @[GameUtilities.scala 21:24]
  reg  _T_363_1; // @[GameUtilities.scala 21:24]
  reg  _T_364_0; // @[GameUtilities.scala 21:24]
  reg  _T_364_1; // @[GameUtilities.scala 21:24]
  wire  _T_365 = _T_363_0 & _T_364_0; // @[SpriteBlender.scala 40:43]
  wire  _T_367 = ~io_datareader_45[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_371_0; // @[GameUtilities.scala 21:24]
  reg  _T_371_1; // @[GameUtilities.scala 21:24]
  reg  _T_372_0; // @[GameUtilities.scala 21:24]
  reg  _T_372_1; // @[GameUtilities.scala 21:24]
  wire  _T_373 = _T_371_0 & _T_372_0; // @[SpriteBlender.scala 40:43]
  wire  _T_375 = ~io_datareader_46[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_379_0; // @[GameUtilities.scala 21:24]
  reg  _T_379_1; // @[GameUtilities.scala 21:24]
  reg  _T_380_0; // @[GameUtilities.scala 21:24]
  reg  _T_380_1; // @[GameUtilities.scala 21:24]
  wire  _T_381 = _T_379_0 & _T_380_0; // @[SpriteBlender.scala 40:43]
  wire  _T_383 = ~io_datareader_47[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_387_0; // @[GameUtilities.scala 21:24]
  reg  _T_387_1; // @[GameUtilities.scala 21:24]
  reg  _T_388_0; // @[GameUtilities.scala 21:24]
  reg  _T_388_1; // @[GameUtilities.scala 21:24]
  wire  _T_389 = _T_387_0 & _T_388_0; // @[SpriteBlender.scala 40:43]
  wire  _T_391 = ~io_datareader_48[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_395_0; // @[GameUtilities.scala 21:24]
  reg  _T_395_1; // @[GameUtilities.scala 21:24]
  reg  _T_396_0; // @[GameUtilities.scala 21:24]
  reg  _T_396_1; // @[GameUtilities.scala 21:24]
  wire  _T_397 = _T_395_0 & _T_396_0; // @[SpriteBlender.scala 40:43]
  wire  _T_399 = ~io_datareader_49[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_403_0; // @[GameUtilities.scala 21:24]
  reg  _T_403_1; // @[GameUtilities.scala 21:24]
  reg  _T_404_0; // @[GameUtilities.scala 21:24]
  reg  _T_404_1; // @[GameUtilities.scala 21:24]
  wire  _T_405 = _T_403_0 & _T_404_0; // @[SpriteBlender.scala 40:43]
  wire  _T_407 = ~io_datareader_50[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_411_0; // @[GameUtilities.scala 21:24]
  reg  _T_411_1; // @[GameUtilities.scala 21:24]
  reg  _T_412_0; // @[GameUtilities.scala 21:24]
  reg  _T_412_1; // @[GameUtilities.scala 21:24]
  wire  _T_413 = _T_411_0 & _T_412_0; // @[SpriteBlender.scala 40:43]
  wire  _T_415 = ~io_datareader_51[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_420_0; // @[GameUtilities.scala 21:24]
  reg  _T_420_1; // @[GameUtilities.scala 21:24]
  wire  _T_423 = ~io_datareader_52[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_428_0; // @[GameUtilities.scala 21:24]
  reg  _T_428_1; // @[GameUtilities.scala 21:24]
  wire  _T_431 = ~io_datareader_53[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_436_0; // @[GameUtilities.scala 21:24]
  reg  _T_436_1; // @[GameUtilities.scala 21:24]
  wire  _T_439 = ~io_datareader_54[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_443_0; // @[GameUtilities.scala 21:24]
  reg  _T_443_1; // @[GameUtilities.scala 21:24]
  reg  _T_444_0; // @[GameUtilities.scala 21:24]
  reg  _T_444_1; // @[GameUtilities.scala 21:24]
  wire  _T_445 = _T_443_0 & _T_444_0; // @[SpriteBlender.scala 40:43]
  wire  _T_447 = ~io_datareader_55[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_451_0; // @[GameUtilities.scala 21:24]
  reg  _T_451_1; // @[GameUtilities.scala 21:24]
  reg  _T_452_0; // @[GameUtilities.scala 21:24]
  reg  _T_452_1; // @[GameUtilities.scala 21:24]
  wire  _T_453 = _T_451_0 & _T_452_0; // @[SpriteBlender.scala 40:43]
  wire  _T_455 = ~io_datareader_56[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_459_0; // @[GameUtilities.scala 21:24]
  reg  _T_459_1; // @[GameUtilities.scala 21:24]
  reg  _T_460_0; // @[GameUtilities.scala 21:24]
  reg  _T_460_1; // @[GameUtilities.scala 21:24]
  wire  _T_461 = _T_459_0 & _T_460_0; // @[SpriteBlender.scala 40:43]
  wire  _T_463 = ~io_datareader_57[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_468_0; // @[GameUtilities.scala 21:24]
  reg  _T_468_1; // @[GameUtilities.scala 21:24]
  wire  _T_471 = ~io_datareader_58[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_476_0; // @[GameUtilities.scala 21:24]
  reg  _T_476_1; // @[GameUtilities.scala 21:24]
  wire  _T_479 = ~io_datareader_59[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_484_0; // @[GameUtilities.scala 21:24]
  reg  _T_484_1; // @[GameUtilities.scala 21:24]
  wire  _T_487 = ~io_datareader_60[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_491_0; // @[GameUtilities.scala 21:24]
  reg  _T_491_1; // @[GameUtilities.scala 21:24]
  reg  _T_492_0; // @[GameUtilities.scala 21:24]
  reg  _T_492_1; // @[GameUtilities.scala 21:24]
  wire  _T_493 = _T_491_0 & _T_492_0; // @[SpriteBlender.scala 40:43]
  wire  _T_495 = ~io_datareader_61[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_499_0; // @[GameUtilities.scala 21:24]
  reg  _T_499_1; // @[GameUtilities.scala 21:24]
  reg  _T_500_0; // @[GameUtilities.scala 21:24]
  reg  _T_500_1; // @[GameUtilities.scala 21:24]
  wire  _T_501 = _T_499_0 & _T_500_0; // @[SpriteBlender.scala 40:43]
  wire  _T_503 = ~io_datareader_62[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_507_0; // @[GameUtilities.scala 21:24]
  reg  _T_507_1; // @[GameUtilities.scala 21:24]
  reg  _T_508_0; // @[GameUtilities.scala 21:24]
  reg  _T_508_1; // @[GameUtilities.scala 21:24]
  wire  _T_509 = _T_507_0 & _T_508_0; // @[SpriteBlender.scala 40:43]
  wire  _T_511 = ~io_datareader_63[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_515_0; // @[GameUtilities.scala 21:24]
  reg  _T_515_1; // @[GameUtilities.scala 21:24]
  reg  _T_516_0; // @[GameUtilities.scala 21:24]
  reg  _T_516_1; // @[GameUtilities.scala 21:24]
  wire  _T_517 = _T_515_0 & _T_516_0; // @[SpriteBlender.scala 40:43]
  wire  _T_519 = ~io_datareader_64[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_523_0; // @[GameUtilities.scala 21:24]
  reg  _T_523_1; // @[GameUtilities.scala 21:24]
  reg  _T_524_0; // @[GameUtilities.scala 21:24]
  reg  _T_524_1; // @[GameUtilities.scala 21:24]
  wire  _T_525 = _T_523_0 & _T_524_0; // @[SpriteBlender.scala 40:43]
  wire  _T_527 = ~io_datareader_65[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_531_0; // @[GameUtilities.scala 21:24]
  reg  _T_531_1; // @[GameUtilities.scala 21:24]
  reg  _T_532_0; // @[GameUtilities.scala 21:24]
  reg  _T_532_1; // @[GameUtilities.scala 21:24]
  wire  _T_533 = _T_531_0 & _T_532_0; // @[SpriteBlender.scala 40:43]
  wire  _T_535 = ~io_datareader_66[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_540_0; // @[GameUtilities.scala 21:24]
  reg  _T_540_1; // @[GameUtilities.scala 21:24]
  wire  _T_543 = ~io_datareader_67[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_548_0; // @[GameUtilities.scala 21:24]
  reg  _T_548_1; // @[GameUtilities.scala 21:24]
  wire  _T_551 = ~io_datareader_68[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_556_0; // @[GameUtilities.scala 21:24]
  reg  _T_556_1; // @[GameUtilities.scala 21:24]
  wire  _T_559 = ~io_datareader_69[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_563_0; // @[GameUtilities.scala 21:24]
  reg  _T_563_1; // @[GameUtilities.scala 21:24]
  reg  _T_564_0; // @[GameUtilities.scala 21:24]
  reg  _T_564_1; // @[GameUtilities.scala 21:24]
  wire  _T_565 = _T_563_0 & _T_564_0; // @[SpriteBlender.scala 40:43]
  wire  _T_567 = ~io_datareader_70[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_571_0; // @[GameUtilities.scala 21:24]
  reg  _T_571_1; // @[GameUtilities.scala 21:24]
  reg  _T_572_0; // @[GameUtilities.scala 21:24]
  reg  _T_572_1; // @[GameUtilities.scala 21:24]
  wire  _T_573 = _T_571_0 & _T_572_0; // @[SpriteBlender.scala 40:43]
  wire  _T_575 = ~io_datareader_71[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_579_0; // @[GameUtilities.scala 21:24]
  reg  _T_579_1; // @[GameUtilities.scala 21:24]
  reg  _T_580_0; // @[GameUtilities.scala 21:24]
  reg  _T_580_1; // @[GameUtilities.scala 21:24]
  wire  _T_581 = _T_579_0 & _T_580_0; // @[SpriteBlender.scala 40:43]
  wire  _T_583 = ~io_datareader_72[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_588_0; // @[GameUtilities.scala 21:24]
  reg  _T_588_1; // @[GameUtilities.scala 21:24]
  wire  _T_591 = ~io_datareader_73[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_596_0; // @[GameUtilities.scala 21:24]
  reg  _T_596_1; // @[GameUtilities.scala 21:24]
  wire  _T_599 = ~io_datareader_74[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_604_0; // @[GameUtilities.scala 21:24]
  reg  _T_604_1; // @[GameUtilities.scala 21:24]
  wire  _T_607 = ~io_datareader_75[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_612_0; // @[GameUtilities.scala 21:24]
  reg  _T_612_1; // @[GameUtilities.scala 21:24]
  wire  _T_615 = ~io_datareader_76[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_620_0; // @[GameUtilities.scala 21:24]
  reg  _T_620_1; // @[GameUtilities.scala 21:24]
  wire  _T_623 = ~io_datareader_77[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_628_0; // @[GameUtilities.scala 21:24]
  reg  _T_628_1; // @[GameUtilities.scala 21:24]
  wire  _T_631 = ~io_datareader_78[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_636_0; // @[GameUtilities.scala 21:24]
  reg  _T_636_1; // @[GameUtilities.scala 21:24]
  wire  _T_639 = ~io_datareader_79[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_644_0; // @[GameUtilities.scala 21:24]
  reg  _T_644_1; // @[GameUtilities.scala 21:24]
  wire  _T_647 = ~io_datareader_80[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_652_0; // @[GameUtilities.scala 21:24]
  reg  _T_652_1; // @[GameUtilities.scala 21:24]
  wire  _T_655 = ~io_datareader_81[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_660_0; // @[GameUtilities.scala 21:24]
  reg  _T_660_1; // @[GameUtilities.scala 21:24]
  wire  _T_663 = ~io_datareader_82[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_668_0; // @[GameUtilities.scala 21:24]
  reg  _T_668_1; // @[GameUtilities.scala 21:24]
  wire  _T_671 = ~io_datareader_83[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_676_0; // @[GameUtilities.scala 21:24]
  reg  _T_676_1; // @[GameUtilities.scala 21:24]
  wire  _T_679 = ~io_datareader_84[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_684_0; // @[GameUtilities.scala 21:24]
  reg  _T_684_1; // @[GameUtilities.scala 21:24]
  wire  _T_687 = ~io_datareader_85[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_692_0; // @[GameUtilities.scala 21:24]
  reg  _T_692_1; // @[GameUtilities.scala 21:24]
  wire  _T_695 = ~io_datareader_86[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_700_0; // @[GameUtilities.scala 21:24]
  reg  _T_700_1; // @[GameUtilities.scala 21:24]
  wire  _T_703 = ~io_datareader_87[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_708_0; // @[GameUtilities.scala 21:24]
  reg  _T_708_1; // @[GameUtilities.scala 21:24]
  wire  _T_711 = ~io_datareader_88[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_716_0; // @[GameUtilities.scala 21:24]
  reg  _T_716_1; // @[GameUtilities.scala 21:24]
  wire  _T_719 = ~io_datareader_89[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_724_0; // @[GameUtilities.scala 21:24]
  reg  _T_724_1; // @[GameUtilities.scala 21:24]
  wire  _T_727 = ~io_datareader_90[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_732_0; // @[GameUtilities.scala 21:24]
  reg  _T_732_1; // @[GameUtilities.scala 21:24]
  wire  _T_735 = ~io_datareader_91[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_740_0; // @[GameUtilities.scala 21:24]
  reg  _T_740_1; // @[GameUtilities.scala 21:24]
  wire  _T_743 = ~io_datareader_92[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_748_0; // @[GameUtilities.scala 21:24]
  reg  _T_748_1; // @[GameUtilities.scala 21:24]
  wire  _T_751 = ~io_datareader_93[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_756_0; // @[GameUtilities.scala 21:24]
  reg  _T_756_1; // @[GameUtilities.scala 21:24]
  wire  _T_759 = ~io_datareader_94[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_764_0; // @[GameUtilities.scala 21:24]
  reg  _T_764_1; // @[GameUtilities.scala 21:24]
  wire  _T_767 = ~io_datareader_95[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_772_0; // @[GameUtilities.scala 21:24]
  reg  _T_772_1; // @[GameUtilities.scala 21:24]
  wire  _T_775 = ~io_datareader_96[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_780_0; // @[GameUtilities.scala 21:24]
  reg  _T_780_1; // @[GameUtilities.scala 21:24]
  wire  _T_783 = ~io_datareader_97[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_788_0; // @[GameUtilities.scala 21:24]
  reg  _T_788_1; // @[GameUtilities.scala 21:24]
  wire  _T_791 = ~io_datareader_98[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_796_0; // @[GameUtilities.scala 21:24]
  reg  _T_796_1; // @[GameUtilities.scala 21:24]
  wire  _T_799 = ~io_datareader_99[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_804_0; // @[GameUtilities.scala 21:24]
  reg  _T_804_1; // @[GameUtilities.scala 21:24]
  wire  _T_807 = ~io_datareader_100[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_812_0; // @[GameUtilities.scala 21:24]
  reg  _T_812_1; // @[GameUtilities.scala 21:24]
  wire  _T_815 = ~io_datareader_101[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_820_0; // @[GameUtilities.scala 21:24]
  reg  _T_820_1; // @[GameUtilities.scala 21:24]
  wire  _T_823 = ~io_datareader_102[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_828_0; // @[GameUtilities.scala 21:24]
  reg  _T_828_1; // @[GameUtilities.scala 21:24]
  wire  _T_831 = ~io_datareader_103[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_836_0; // @[GameUtilities.scala 21:24]
  reg  _T_836_1; // @[GameUtilities.scala 21:24]
  wire  _T_839 = ~io_datareader_104[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_844_0; // @[GameUtilities.scala 21:24]
  reg  _T_844_1; // @[GameUtilities.scala 21:24]
  wire  _T_847 = ~io_datareader_105[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_852_0; // @[GameUtilities.scala 21:24]
  reg  _T_852_1; // @[GameUtilities.scala 21:24]
  wire  _T_855 = ~io_datareader_106[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_860_0; // @[GameUtilities.scala 21:24]
  reg  _T_860_1; // @[GameUtilities.scala 21:24]
  wire  _T_863 = ~io_datareader_107[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_868_0; // @[GameUtilities.scala 21:24]
  reg  _T_868_1; // @[GameUtilities.scala 21:24]
  wire  _T_871 = ~io_datareader_108[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_876_0; // @[GameUtilities.scala 21:24]
  reg  _T_876_1; // @[GameUtilities.scala 21:24]
  wire  _T_879 = ~io_datareader_109[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_884_0; // @[GameUtilities.scala 21:24]
  reg  _T_884_1; // @[GameUtilities.scala 21:24]
  wire  _T_887 = ~io_datareader_110[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_892_0; // @[GameUtilities.scala 21:24]
  reg  _T_892_1; // @[GameUtilities.scala 21:24]
  wire  _T_895 = ~io_datareader_111[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_900_0; // @[GameUtilities.scala 21:24]
  reg  _T_900_1; // @[GameUtilities.scala 21:24]
  wire  _T_903 = ~io_datareader_112[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_908_0; // @[GameUtilities.scala 21:24]
  reg  _T_908_1; // @[GameUtilities.scala 21:24]
  wire  _T_911 = ~io_datareader_113[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_916_0; // @[GameUtilities.scala 21:24]
  reg  _T_916_1; // @[GameUtilities.scala 21:24]
  wire  _T_919 = ~io_datareader_114[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_924_0; // @[GameUtilities.scala 21:24]
  reg  _T_924_1; // @[GameUtilities.scala 21:24]
  wire  _T_927 = ~io_datareader_115[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_932_0; // @[GameUtilities.scala 21:24]
  reg  _T_932_1; // @[GameUtilities.scala 21:24]
  wire  _T_935 = ~io_datareader_116[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_940_0; // @[GameUtilities.scala 21:24]
  reg  _T_940_1; // @[GameUtilities.scala 21:24]
  wire  _T_943 = ~io_datareader_117[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_948_0; // @[GameUtilities.scala 21:24]
  reg  _T_948_1; // @[GameUtilities.scala 21:24]
  wire  _T_951 = ~io_datareader_118[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_956_0; // @[GameUtilities.scala 21:24]
  reg  _T_956_1; // @[GameUtilities.scala 21:24]
  wire  _T_959 = ~io_datareader_119[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_964_0; // @[GameUtilities.scala 21:24]
  reg  _T_964_1; // @[GameUtilities.scala 21:24]
  wire  _T_967 = ~io_datareader_120[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_972_0; // @[GameUtilities.scala 21:24]
  reg  _T_972_1; // @[GameUtilities.scala 21:24]
  wire  _T_975 = ~io_datareader_121[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_980_0; // @[GameUtilities.scala 21:24]
  reg  _T_980_1; // @[GameUtilities.scala 21:24]
  wire  _T_983 = ~io_datareader_122[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_988_0; // @[GameUtilities.scala 21:24]
  reg  _T_988_1; // @[GameUtilities.scala 21:24]
  wire  _T_991 = ~io_datareader_123[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_996_0; // @[GameUtilities.scala 21:24]
  reg  _T_996_1; // @[GameUtilities.scala 21:24]
  wire  _T_999 = ~io_datareader_124[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_1004_0; // @[GameUtilities.scala 21:24]
  reg  _T_1004_1; // @[GameUtilities.scala 21:24]
  wire  _T_1007 = ~io_datareader_125[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_1012_0; // @[GameUtilities.scala 21:24]
  reg  _T_1012_1; // @[GameUtilities.scala 21:24]
  wire  _T_1015 = ~io_datareader_126[6]; // @[SpriteBlender.scala 42:9]
  reg  _T_1020_0; // @[GameUtilities.scala 21:24]
  reg  _T_1020_1; // @[GameUtilities.scala 21:24]
  wire  _T_1023 = ~io_datareader_127[6]; // @[SpriteBlender.scala 42:9]
  wire  topSpriteAlpha = multiHotPriortyReductionTree_io_dataOutput[6]; // @[SpriteBlender.scala 49:38]
  wire [5:0] topSpriteRGB = multiHotPriortyReductionTree_io_dataOutput[5:0]; // @[SpriteBlender.scala 50:36]
  reg  _T_1026_0; // @[GameUtilities.scala 21:24]
  reg  _T_1026_1; // @[GameUtilities.scala 21:24]
  reg  _T_1027_0; // @[GameUtilities.scala 21:24]
  reg  _T_1027_1; // @[GameUtilities.scala 21:24]
  wire  _T_1029 = _T_1026_0 & _T_1027_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1032 = _T_1029 & _T_7; // @[SpriteBlender.scala 63:35]
  wire  _T_1033 = 7'h0 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_0 = _T_1032 & _T_1033; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_0 = io_datareader_0[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1038_0; // @[GameUtilities.scala 21:24]
  reg  _T_1038_1; // @[GameUtilities.scala 21:24]
  reg  _T_1039_0; // @[GameUtilities.scala 21:24]
  reg  _T_1039_1; // @[GameUtilities.scala 21:24]
  wire  _T_1041 = _T_1038_0 & _T_1039_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1044 = _T_1041 & _T_15; // @[SpriteBlender.scala 63:35]
  wire  _T_1045 = 7'h1 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_1 = _T_1044 & _T_1045; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_1 = io_datareader_1[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1050_0; // @[GameUtilities.scala 21:24]
  reg  _T_1050_1; // @[GameUtilities.scala 21:24]
  reg  _T_1051_0; // @[GameUtilities.scala 21:24]
  reg  _T_1051_1; // @[GameUtilities.scala 21:24]
  wire  _T_1053 = _T_1050_0 & _T_1051_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1056 = _T_1053 & _T_23; // @[SpriteBlender.scala 63:35]
  wire  _T_1057 = 7'h2 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_2 = _T_1056 & _T_1057; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_2 = io_datareader_2[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1062_0; // @[GameUtilities.scala 21:24]
  reg  _T_1062_1; // @[GameUtilities.scala 21:24]
  reg  _T_1063_0; // @[GameUtilities.scala 21:24]
  reg  _T_1063_1; // @[GameUtilities.scala 21:24]
  wire  _T_1065 = _T_1062_0 & _T_1063_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1068 = _T_1065 & _T_31; // @[SpriteBlender.scala 63:35]
  wire  _T_1069 = 7'h3 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_3 = _T_1068 & _T_1069; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_3 = io_datareader_3[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1074_0; // @[GameUtilities.scala 21:24]
  reg  _T_1074_1; // @[GameUtilities.scala 21:24]
  reg  _T_1075_0; // @[GameUtilities.scala 21:24]
  reg  _T_1075_1; // @[GameUtilities.scala 21:24]
  wire  _T_1077 = _T_1074_0 & _T_1075_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1080 = _T_1077 & _T_39; // @[SpriteBlender.scala 63:35]
  wire  _T_1081 = 7'h4 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_4 = _T_1080 & _T_1081; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_4 = io_datareader_4[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1086_0; // @[GameUtilities.scala 21:24]
  reg  _T_1086_1; // @[GameUtilities.scala 21:24]
  reg  _T_1087_0; // @[GameUtilities.scala 21:24]
  reg  _T_1087_1; // @[GameUtilities.scala 21:24]
  wire  _T_1089 = _T_1086_0 & _T_1087_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1092 = _T_1089 & _T_47; // @[SpriteBlender.scala 63:35]
  wire  _T_1093 = 7'h5 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_5 = _T_1092 & _T_1093; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_5 = io_datareader_5[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1098_0; // @[GameUtilities.scala 21:24]
  reg  _T_1098_1; // @[GameUtilities.scala 21:24]
  reg  _T_1099_0; // @[GameUtilities.scala 21:24]
  reg  _T_1099_1; // @[GameUtilities.scala 21:24]
  wire  _T_1101 = _T_1098_0 & _T_1099_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1104 = _T_1101 & _T_55; // @[SpriteBlender.scala 63:35]
  wire  _T_1105 = 7'h6 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_6 = _T_1104 & _T_1105; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_6 = io_datareader_6[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1110_0; // @[GameUtilities.scala 21:24]
  reg  _T_1110_1; // @[GameUtilities.scala 21:24]
  reg  _T_1111_0; // @[GameUtilities.scala 21:24]
  reg  _T_1111_1; // @[GameUtilities.scala 21:24]
  wire  _T_1113 = _T_1110_0 & _T_1111_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1116 = _T_1113 & _T_63; // @[SpriteBlender.scala 63:35]
  wire  _T_1117 = 7'h7 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_7 = _T_1116 & _T_1117; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_7 = io_datareader_7[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1122_0; // @[GameUtilities.scala 21:24]
  reg  _T_1122_1; // @[GameUtilities.scala 21:24]
  reg  _T_1123_0; // @[GameUtilities.scala 21:24]
  reg  _T_1123_1; // @[GameUtilities.scala 21:24]
  wire  _T_1125 = _T_1122_0 & _T_1123_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1128 = _T_1125 & _T_71; // @[SpriteBlender.scala 63:35]
  wire  _T_1129 = 7'h8 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_8 = _T_1128 & _T_1129; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_8 = io_datareader_8[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1134_0; // @[GameUtilities.scala 21:24]
  reg  _T_1134_1; // @[GameUtilities.scala 21:24]
  reg  _T_1135_0; // @[GameUtilities.scala 21:24]
  reg  _T_1135_1; // @[GameUtilities.scala 21:24]
  wire  _T_1137 = _T_1134_0 & _T_1135_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1140 = _T_1137 & _T_79; // @[SpriteBlender.scala 63:35]
  wire  _T_1141 = 7'h9 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_9 = _T_1140 & _T_1141; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_9 = io_datareader_9[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1146_0; // @[GameUtilities.scala 21:24]
  reg  _T_1146_1; // @[GameUtilities.scala 21:24]
  reg  _T_1147_0; // @[GameUtilities.scala 21:24]
  reg  _T_1147_1; // @[GameUtilities.scala 21:24]
  wire  _T_1149 = _T_1146_0 & _T_1147_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1152 = _T_1149 & _T_87; // @[SpriteBlender.scala 63:35]
  wire  _T_1153 = 7'ha != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_10 = _T_1152 & _T_1153; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_10 = io_datareader_10[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1158_0; // @[GameUtilities.scala 21:24]
  reg  _T_1158_1; // @[GameUtilities.scala 21:24]
  reg  _T_1159_0; // @[GameUtilities.scala 21:24]
  reg  _T_1159_1; // @[GameUtilities.scala 21:24]
  wire  _T_1161 = _T_1158_0 & _T_1159_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1164 = _T_1161 & _T_95; // @[SpriteBlender.scala 63:35]
  wire  _T_1165 = 7'hb != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_11 = _T_1164 & _T_1165; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_11 = io_datareader_11[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1170_0; // @[GameUtilities.scala 21:24]
  reg  _T_1170_1; // @[GameUtilities.scala 21:24]
  reg  _T_1171_0; // @[GameUtilities.scala 21:24]
  reg  _T_1171_1; // @[GameUtilities.scala 21:24]
  wire  _T_1173 = _T_1170_0 & _T_1171_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1176 = _T_1173 & _T_103; // @[SpriteBlender.scala 63:35]
  wire  _T_1177 = 7'hc != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_12 = _T_1176 & _T_1177; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_12 = io_datareader_12[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1182_0; // @[GameUtilities.scala 21:24]
  reg  _T_1182_1; // @[GameUtilities.scala 21:24]
  reg  _T_1183_0; // @[GameUtilities.scala 21:24]
  reg  _T_1183_1; // @[GameUtilities.scala 21:24]
  wire  _T_1185 = _T_1182_0 & _T_1183_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1188 = _T_1185 & _T_111; // @[SpriteBlender.scala 63:35]
  wire  _T_1189 = 7'hd != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_13 = _T_1188 & _T_1189; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_13 = io_datareader_13[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1194_0; // @[GameUtilities.scala 21:24]
  reg  _T_1194_1; // @[GameUtilities.scala 21:24]
  reg  _T_1195_0; // @[GameUtilities.scala 21:24]
  reg  _T_1195_1; // @[GameUtilities.scala 21:24]
  wire  _T_1197 = _T_1194_0 & _T_1195_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1200 = _T_1197 & _T_119; // @[SpriteBlender.scala 63:35]
  wire  _T_1201 = 7'he != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_14 = _T_1200 & _T_1201; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_14 = io_datareader_14[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1206_0; // @[GameUtilities.scala 21:24]
  reg  _T_1206_1; // @[GameUtilities.scala 21:24]
  reg  _T_1207_0; // @[GameUtilities.scala 21:24]
  reg  _T_1207_1; // @[GameUtilities.scala 21:24]
  wire  _T_1209 = _T_1206_0 & _T_1207_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1212 = _T_1209 & _T_127; // @[SpriteBlender.scala 63:35]
  wire  _T_1213 = 7'hf != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_15 = _T_1212 & _T_1213; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_15 = io_datareader_15[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1218_0; // @[GameUtilities.scala 21:24]
  reg  _T_1218_1; // @[GameUtilities.scala 21:24]
  reg  _T_1219_0; // @[GameUtilities.scala 21:24]
  reg  _T_1219_1; // @[GameUtilities.scala 21:24]
  wire  _T_1221 = _T_1218_0 & _T_1219_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1224 = _T_1221 & _T_135; // @[SpriteBlender.scala 63:35]
  wire  _T_1225 = 7'h10 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_16 = _T_1224 & _T_1225; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_16 = io_datareader_16[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1230_0; // @[GameUtilities.scala 21:24]
  reg  _T_1230_1; // @[GameUtilities.scala 21:24]
  reg  _T_1231_0; // @[GameUtilities.scala 21:24]
  reg  _T_1231_1; // @[GameUtilities.scala 21:24]
  wire  _T_1233 = _T_1230_0 & _T_1231_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1236 = _T_1233 & _T_143; // @[SpriteBlender.scala 63:35]
  wire  _T_1237 = 7'h11 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_17 = _T_1236 & _T_1237; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_17 = io_datareader_17[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1242_0; // @[GameUtilities.scala 21:24]
  reg  _T_1242_1; // @[GameUtilities.scala 21:24]
  reg  _T_1243_0; // @[GameUtilities.scala 21:24]
  reg  _T_1243_1; // @[GameUtilities.scala 21:24]
  wire  _T_1245 = _T_1242_0 & _T_1243_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1248 = _T_1245 & _T_151; // @[SpriteBlender.scala 63:35]
  wire  _T_1249 = 7'h12 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_18 = _T_1248 & _T_1249; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_18 = io_datareader_18[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1254_0; // @[GameUtilities.scala 21:24]
  reg  _T_1254_1; // @[GameUtilities.scala 21:24]
  reg  _T_1255_0; // @[GameUtilities.scala 21:24]
  reg  _T_1255_1; // @[GameUtilities.scala 21:24]
  wire  _T_1257 = _T_1254_0 & _T_1255_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1260 = _T_1257 & _T_159; // @[SpriteBlender.scala 63:35]
  wire  _T_1261 = 7'h13 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_19 = _T_1260 & _T_1261; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_19 = io_datareader_19[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1266_0; // @[GameUtilities.scala 21:24]
  reg  _T_1266_1; // @[GameUtilities.scala 21:24]
  reg  _T_1267_0; // @[GameUtilities.scala 21:24]
  reg  _T_1267_1; // @[GameUtilities.scala 21:24]
  wire  _T_1269 = _T_1266_0 & _T_1267_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1272 = _T_1269 & _T_167; // @[SpriteBlender.scala 63:35]
  wire  _T_1273 = 7'h14 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_20 = _T_1272 & _T_1273; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_20 = io_datareader_20[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1278_0; // @[GameUtilities.scala 21:24]
  reg  _T_1278_1; // @[GameUtilities.scala 21:24]
  reg  _T_1279_0; // @[GameUtilities.scala 21:24]
  reg  _T_1279_1; // @[GameUtilities.scala 21:24]
  wire  _T_1281 = _T_1278_0 & _T_1279_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1284 = _T_1281 & _T_175; // @[SpriteBlender.scala 63:35]
  wire  _T_1285 = 7'h15 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_21 = _T_1284 & _T_1285; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_21 = io_datareader_21[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1290_0; // @[GameUtilities.scala 21:24]
  reg  _T_1290_1; // @[GameUtilities.scala 21:24]
  reg  _T_1291_0; // @[GameUtilities.scala 21:24]
  reg  _T_1291_1; // @[GameUtilities.scala 21:24]
  wire  _T_1293 = _T_1290_0 & _T_1291_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1296 = _T_1293 & _T_183; // @[SpriteBlender.scala 63:35]
  wire  _T_1297 = 7'h16 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_22 = _T_1296 & _T_1297; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_22 = io_datareader_22[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1302_0; // @[GameUtilities.scala 21:24]
  reg  _T_1302_1; // @[GameUtilities.scala 21:24]
  reg  _T_1303_0; // @[GameUtilities.scala 21:24]
  reg  _T_1303_1; // @[GameUtilities.scala 21:24]
  wire  _T_1305 = _T_1302_0 & _T_1303_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1308 = _T_1305 & _T_191; // @[SpriteBlender.scala 63:35]
  wire  _T_1309 = 7'h17 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_23 = _T_1308 & _T_1309; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_23 = io_datareader_23[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1314_0; // @[GameUtilities.scala 21:24]
  reg  _T_1314_1; // @[GameUtilities.scala 21:24]
  reg  _T_1315_0; // @[GameUtilities.scala 21:24]
  reg  _T_1315_1; // @[GameUtilities.scala 21:24]
  wire  _T_1317 = _T_1314_0 & _T_1315_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1320 = _T_1317 & _T_199; // @[SpriteBlender.scala 63:35]
  wire  _T_1321 = 7'h18 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_24 = _T_1320 & _T_1321; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_24 = io_datareader_24[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1326_0; // @[GameUtilities.scala 21:24]
  reg  _T_1326_1; // @[GameUtilities.scala 21:24]
  reg  _T_1327_0; // @[GameUtilities.scala 21:24]
  reg  _T_1327_1; // @[GameUtilities.scala 21:24]
  wire  _T_1329 = _T_1326_0 & _T_1327_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1332 = _T_1329 & _T_207; // @[SpriteBlender.scala 63:35]
  wire  _T_1333 = 7'h19 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_25 = _T_1332 & _T_1333; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_25 = io_datareader_25[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1338_0; // @[GameUtilities.scala 21:24]
  reg  _T_1338_1; // @[GameUtilities.scala 21:24]
  reg  _T_1339_0; // @[GameUtilities.scala 21:24]
  reg  _T_1339_1; // @[GameUtilities.scala 21:24]
  wire  _T_1341 = _T_1338_0 & _T_1339_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1344 = _T_1341 & _T_215; // @[SpriteBlender.scala 63:35]
  wire  _T_1345 = 7'h1a != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_26 = _T_1344 & _T_1345; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_26 = io_datareader_26[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1350_0; // @[GameUtilities.scala 21:24]
  reg  _T_1350_1; // @[GameUtilities.scala 21:24]
  reg  _T_1351_0; // @[GameUtilities.scala 21:24]
  reg  _T_1351_1; // @[GameUtilities.scala 21:24]
  wire  _T_1353 = _T_1350_0 & _T_1351_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1356 = _T_1353 & _T_223; // @[SpriteBlender.scala 63:35]
  wire  _T_1357 = 7'h1b != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_27 = _T_1356 & _T_1357; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_27 = io_datareader_27[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1362_0; // @[GameUtilities.scala 21:24]
  reg  _T_1362_1; // @[GameUtilities.scala 21:24]
  reg  _T_1363_0; // @[GameUtilities.scala 21:24]
  reg  _T_1363_1; // @[GameUtilities.scala 21:24]
  wire  _T_1365 = _T_1362_0 & _T_1363_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1368 = _T_1365 & _T_231; // @[SpriteBlender.scala 63:35]
  wire  _T_1369 = 7'h1c != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_28 = _T_1368 & _T_1369; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_28 = io_datareader_28[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1374_0; // @[GameUtilities.scala 21:24]
  reg  _T_1374_1; // @[GameUtilities.scala 21:24]
  reg  _T_1375_0; // @[GameUtilities.scala 21:24]
  reg  _T_1375_1; // @[GameUtilities.scala 21:24]
  wire  _T_1377 = _T_1374_0 & _T_1375_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1380 = _T_1377 & _T_239; // @[SpriteBlender.scala 63:35]
  wire  _T_1381 = 7'h1d != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_29 = _T_1380 & _T_1381; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_29 = io_datareader_29[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1386_0; // @[GameUtilities.scala 21:24]
  reg  _T_1386_1; // @[GameUtilities.scala 21:24]
  reg  _T_1387_0; // @[GameUtilities.scala 21:24]
  reg  _T_1387_1; // @[GameUtilities.scala 21:24]
  wire  _T_1389 = _T_1386_0 & _T_1387_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1392 = _T_1389 & _T_247; // @[SpriteBlender.scala 63:35]
  wire  _T_1393 = 7'h1e != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_30 = _T_1392 & _T_1393; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_30 = io_datareader_30[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1398_0; // @[GameUtilities.scala 21:24]
  reg  _T_1398_1; // @[GameUtilities.scala 21:24]
  reg  _T_1399_0; // @[GameUtilities.scala 21:24]
  reg  _T_1399_1; // @[GameUtilities.scala 21:24]
  wire  _T_1401 = _T_1398_0 & _T_1399_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1404 = _T_1401 & _T_255; // @[SpriteBlender.scala 63:35]
  wire  _T_1405 = 7'h1f != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_31 = _T_1404 & _T_1405; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_31 = io_datareader_31[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1410_0; // @[GameUtilities.scala 21:24]
  reg  _T_1410_1; // @[GameUtilities.scala 21:24]
  reg  _T_1411_0; // @[GameUtilities.scala 21:24]
  reg  _T_1411_1; // @[GameUtilities.scala 21:24]
  wire  _T_1413 = _T_1410_0 & _T_1411_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1416 = _T_1413 & _T_263; // @[SpriteBlender.scala 63:35]
  wire  _T_1417 = 7'h20 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_32 = _T_1416 & _T_1417; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_32 = io_datareader_32[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1422_0; // @[GameUtilities.scala 21:24]
  reg  _T_1422_1; // @[GameUtilities.scala 21:24]
  reg  _T_1423_0; // @[GameUtilities.scala 21:24]
  reg  _T_1423_1; // @[GameUtilities.scala 21:24]
  wire  _T_1425 = _T_1422_0 & _T_1423_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1428 = _T_1425 & _T_271; // @[SpriteBlender.scala 63:35]
  wire  _T_1429 = 7'h21 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_33 = _T_1428 & _T_1429; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_33 = io_datareader_33[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1435_0; // @[GameUtilities.scala 21:24]
  reg  _T_1435_1; // @[GameUtilities.scala 21:24]
  wire  _T_1440 = _T_1435_0 & _T_279; // @[SpriteBlender.scala 63:35]
  wire  _T_1441 = 7'h22 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_34 = _T_1440 & _T_1441; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_34 = io_datareader_34[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1447_0; // @[GameUtilities.scala 21:24]
  reg  _T_1447_1; // @[GameUtilities.scala 21:24]
  wire  _T_1452 = _T_1447_0 & _T_287; // @[SpriteBlender.scala 63:35]
  wire  _T_1453 = 7'h23 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_35 = _T_1452 & _T_1453; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_35 = io_datareader_35[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1459_0; // @[GameUtilities.scala 21:24]
  reg  _T_1459_1; // @[GameUtilities.scala 21:24]
  wire  _T_1464 = _T_1459_0 & _T_295; // @[SpriteBlender.scala 63:35]
  wire  _T_1465 = 7'h24 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_36 = _T_1464 & _T_1465; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_36 = io_datareader_36[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1471_0; // @[GameUtilities.scala 21:24]
  reg  _T_1471_1; // @[GameUtilities.scala 21:24]
  wire  _T_1476 = _T_1471_0 & _T_303; // @[SpriteBlender.scala 63:35]
  wire  _T_1477 = 7'h25 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_37 = _T_1476 & _T_1477; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_37 = io_datareader_37[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1483_0; // @[GameUtilities.scala 21:24]
  reg  _T_1483_1; // @[GameUtilities.scala 21:24]
  wire  _T_1488 = _T_1483_0 & _T_311; // @[SpriteBlender.scala 63:35]
  wire  _T_1489 = 7'h26 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_38 = _T_1488 & _T_1489; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_38 = io_datareader_38[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1495_0; // @[GameUtilities.scala 21:24]
  reg  _T_1495_1; // @[GameUtilities.scala 21:24]
  wire  _T_1500 = _T_1495_0 & _T_319; // @[SpriteBlender.scala 63:35]
  wire  _T_1501 = 7'h27 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_39 = _T_1500 & _T_1501; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_39 = io_datareader_39[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1507_0; // @[GameUtilities.scala 21:24]
  reg  _T_1507_1; // @[GameUtilities.scala 21:24]
  wire  _T_1512 = _T_1507_0 & _T_327; // @[SpriteBlender.scala 63:35]
  wire  _T_1513 = 7'h28 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_40 = _T_1512 & _T_1513; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_40 = io_datareader_40[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1518_0; // @[GameUtilities.scala 21:24]
  reg  _T_1518_1; // @[GameUtilities.scala 21:24]
  reg  _T_1519_0; // @[GameUtilities.scala 21:24]
  reg  _T_1519_1; // @[GameUtilities.scala 21:24]
  wire  _T_1521 = _T_1518_0 & _T_1519_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1524 = _T_1521 & _T_335; // @[SpriteBlender.scala 63:35]
  wire  _T_1525 = 7'h29 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_41 = _T_1524 & _T_1525; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_41 = io_datareader_41[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1530_0; // @[GameUtilities.scala 21:24]
  reg  _T_1530_1; // @[GameUtilities.scala 21:24]
  reg  _T_1531_0; // @[GameUtilities.scala 21:24]
  reg  _T_1531_1; // @[GameUtilities.scala 21:24]
  wire  _T_1533 = _T_1530_0 & _T_1531_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1536 = _T_1533 & _T_343; // @[SpriteBlender.scala 63:35]
  wire  _T_1537 = 7'h2a != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_42 = _T_1536 & _T_1537; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_42 = io_datareader_42[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1542_0; // @[GameUtilities.scala 21:24]
  reg  _T_1542_1; // @[GameUtilities.scala 21:24]
  reg  _T_1543_0; // @[GameUtilities.scala 21:24]
  reg  _T_1543_1; // @[GameUtilities.scala 21:24]
  wire  _T_1545 = _T_1542_0 & _T_1543_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1548 = _T_1545 & _T_351; // @[SpriteBlender.scala 63:35]
  wire  _T_1549 = 7'h2b != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_43 = _T_1548 & _T_1549; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_43 = io_datareader_43[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1554_0; // @[GameUtilities.scala 21:24]
  reg  _T_1554_1; // @[GameUtilities.scala 21:24]
  reg  _T_1555_0; // @[GameUtilities.scala 21:24]
  reg  _T_1555_1; // @[GameUtilities.scala 21:24]
  wire  _T_1557 = _T_1554_0 & _T_1555_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1560 = _T_1557 & _T_359; // @[SpriteBlender.scala 63:35]
  wire  _T_1561 = 7'h2c != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_44 = _T_1560 & _T_1561; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_44 = io_datareader_44[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1566_0; // @[GameUtilities.scala 21:24]
  reg  _T_1566_1; // @[GameUtilities.scala 21:24]
  reg  _T_1567_0; // @[GameUtilities.scala 21:24]
  reg  _T_1567_1; // @[GameUtilities.scala 21:24]
  wire  _T_1569 = _T_1566_0 & _T_1567_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1572 = _T_1569 & _T_367; // @[SpriteBlender.scala 63:35]
  wire  _T_1573 = 7'h2d != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_45 = _T_1572 & _T_1573; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_45 = io_datareader_45[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1578_0; // @[GameUtilities.scala 21:24]
  reg  _T_1578_1; // @[GameUtilities.scala 21:24]
  reg  _T_1579_0; // @[GameUtilities.scala 21:24]
  reg  _T_1579_1; // @[GameUtilities.scala 21:24]
  wire  _T_1581 = _T_1578_0 & _T_1579_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1584 = _T_1581 & _T_375; // @[SpriteBlender.scala 63:35]
  wire  _T_1585 = 7'h2e != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_46 = _T_1584 & _T_1585; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_46 = io_datareader_46[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1590_0; // @[GameUtilities.scala 21:24]
  reg  _T_1590_1; // @[GameUtilities.scala 21:24]
  reg  _T_1591_0; // @[GameUtilities.scala 21:24]
  reg  _T_1591_1; // @[GameUtilities.scala 21:24]
  wire  _T_1593 = _T_1590_0 & _T_1591_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1596 = _T_1593 & _T_383; // @[SpriteBlender.scala 63:35]
  wire  _T_1597 = 7'h2f != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_47 = _T_1596 & _T_1597; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_47 = io_datareader_47[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1602_0; // @[GameUtilities.scala 21:24]
  reg  _T_1602_1; // @[GameUtilities.scala 21:24]
  reg  _T_1603_0; // @[GameUtilities.scala 21:24]
  reg  _T_1603_1; // @[GameUtilities.scala 21:24]
  wire  _T_1605 = _T_1602_0 & _T_1603_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1608 = _T_1605 & _T_391; // @[SpriteBlender.scala 63:35]
  wire  _T_1609 = 7'h30 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_48 = _T_1608 & _T_1609; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_48 = io_datareader_48[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1614_0; // @[GameUtilities.scala 21:24]
  reg  _T_1614_1; // @[GameUtilities.scala 21:24]
  reg  _T_1615_0; // @[GameUtilities.scala 21:24]
  reg  _T_1615_1; // @[GameUtilities.scala 21:24]
  wire  _T_1617 = _T_1614_0 & _T_1615_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1620 = _T_1617 & _T_399; // @[SpriteBlender.scala 63:35]
  wire  _T_1621 = 7'h31 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_49 = _T_1620 & _T_1621; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_49 = io_datareader_49[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1626_0; // @[GameUtilities.scala 21:24]
  reg  _T_1626_1; // @[GameUtilities.scala 21:24]
  reg  _T_1627_0; // @[GameUtilities.scala 21:24]
  reg  _T_1627_1; // @[GameUtilities.scala 21:24]
  wire  _T_1629 = _T_1626_0 & _T_1627_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1632 = _T_1629 & _T_407; // @[SpriteBlender.scala 63:35]
  wire  _T_1633 = 7'h32 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_50 = _T_1632 & _T_1633; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_50 = io_datareader_50[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1638_0; // @[GameUtilities.scala 21:24]
  reg  _T_1638_1; // @[GameUtilities.scala 21:24]
  reg  _T_1639_0; // @[GameUtilities.scala 21:24]
  reg  _T_1639_1; // @[GameUtilities.scala 21:24]
  wire  _T_1641 = _T_1638_0 & _T_1639_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1644 = _T_1641 & _T_415; // @[SpriteBlender.scala 63:35]
  wire  _T_1645 = 7'h33 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_51 = _T_1644 & _T_1645; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_51 = io_datareader_51[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1651_0; // @[GameUtilities.scala 21:24]
  reg  _T_1651_1; // @[GameUtilities.scala 21:24]
  wire  _T_1656 = _T_1651_0 & _T_423; // @[SpriteBlender.scala 63:35]
  wire  _T_1657 = 7'h34 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_52 = _T_1656 & _T_1657; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_52 = io_datareader_52[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1663_0; // @[GameUtilities.scala 21:24]
  reg  _T_1663_1; // @[GameUtilities.scala 21:24]
  wire  _T_1668 = _T_1663_0 & _T_431; // @[SpriteBlender.scala 63:35]
  wire  _T_1669 = 7'h35 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_53 = _T_1668 & _T_1669; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_53 = io_datareader_53[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1675_0; // @[GameUtilities.scala 21:24]
  reg  _T_1675_1; // @[GameUtilities.scala 21:24]
  wire  _T_1680 = _T_1675_0 & _T_439; // @[SpriteBlender.scala 63:35]
  wire  _T_1681 = 7'h36 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_54 = _T_1680 & _T_1681; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_54 = io_datareader_54[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1686_0; // @[GameUtilities.scala 21:24]
  reg  _T_1686_1; // @[GameUtilities.scala 21:24]
  reg  _T_1687_0; // @[GameUtilities.scala 21:24]
  reg  _T_1687_1; // @[GameUtilities.scala 21:24]
  wire  _T_1689 = _T_1686_0 & _T_1687_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1692 = _T_1689 & _T_447; // @[SpriteBlender.scala 63:35]
  wire  _T_1693 = 7'h37 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_55 = _T_1692 & _T_1693; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_55 = io_datareader_55[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1698_0; // @[GameUtilities.scala 21:24]
  reg  _T_1698_1; // @[GameUtilities.scala 21:24]
  reg  _T_1699_0; // @[GameUtilities.scala 21:24]
  reg  _T_1699_1; // @[GameUtilities.scala 21:24]
  wire  _T_1701 = _T_1698_0 & _T_1699_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1704 = _T_1701 & _T_455; // @[SpriteBlender.scala 63:35]
  wire  _T_1705 = 7'h38 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_56 = _T_1704 & _T_1705; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_56 = io_datareader_56[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1710_0; // @[GameUtilities.scala 21:24]
  reg  _T_1710_1; // @[GameUtilities.scala 21:24]
  reg  _T_1711_0; // @[GameUtilities.scala 21:24]
  reg  _T_1711_1; // @[GameUtilities.scala 21:24]
  wire  _T_1713 = _T_1710_0 & _T_1711_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1716 = _T_1713 & _T_463; // @[SpriteBlender.scala 63:35]
  wire  _T_1717 = 7'h39 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_57 = _T_1716 & _T_1717; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_57 = io_datareader_57[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1723_0; // @[GameUtilities.scala 21:24]
  reg  _T_1723_1; // @[GameUtilities.scala 21:24]
  wire  _T_1728 = _T_1723_0 & _T_471; // @[SpriteBlender.scala 63:35]
  wire  _T_1729 = 7'h3a != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_58 = _T_1728 & _T_1729; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_58 = io_datareader_58[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1735_0; // @[GameUtilities.scala 21:24]
  reg  _T_1735_1; // @[GameUtilities.scala 21:24]
  wire  _T_1740 = _T_1735_0 & _T_479; // @[SpriteBlender.scala 63:35]
  wire  _T_1741 = 7'h3b != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_59 = _T_1740 & _T_1741; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_59 = io_datareader_59[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1747_0; // @[GameUtilities.scala 21:24]
  reg  _T_1747_1; // @[GameUtilities.scala 21:24]
  wire  _T_1752 = _T_1747_0 & _T_487; // @[SpriteBlender.scala 63:35]
  wire  _T_1753 = 7'h3c != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_60 = _T_1752 & _T_1753; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_60 = io_datareader_60[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1758_0; // @[GameUtilities.scala 21:24]
  reg  _T_1758_1; // @[GameUtilities.scala 21:24]
  reg  _T_1759_0; // @[GameUtilities.scala 21:24]
  reg  _T_1759_1; // @[GameUtilities.scala 21:24]
  wire  _T_1761 = _T_1758_0 & _T_1759_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1764 = _T_1761 & _T_495; // @[SpriteBlender.scala 63:35]
  wire  _T_1765 = 7'h3d != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_61 = _T_1764 & _T_1765; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_61 = io_datareader_61[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1770_0; // @[GameUtilities.scala 21:24]
  reg  _T_1770_1; // @[GameUtilities.scala 21:24]
  reg  _T_1771_0; // @[GameUtilities.scala 21:24]
  reg  _T_1771_1; // @[GameUtilities.scala 21:24]
  wire  _T_1773 = _T_1770_0 & _T_1771_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1776 = _T_1773 & _T_503; // @[SpriteBlender.scala 63:35]
  wire  _T_1777 = 7'h3e != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_62 = _T_1776 & _T_1777; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_62 = io_datareader_62[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1782_0; // @[GameUtilities.scala 21:24]
  reg  _T_1782_1; // @[GameUtilities.scala 21:24]
  reg  _T_1783_0; // @[GameUtilities.scala 21:24]
  reg  _T_1783_1; // @[GameUtilities.scala 21:24]
  wire  _T_1785 = _T_1782_0 & _T_1783_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1788 = _T_1785 & _T_511; // @[SpriteBlender.scala 63:35]
  wire  _T_1789 = 7'h3f != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_63 = _T_1788 & _T_1789; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_63 = io_datareader_63[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1794_0; // @[GameUtilities.scala 21:24]
  reg  _T_1794_1; // @[GameUtilities.scala 21:24]
  reg  _T_1795_0; // @[GameUtilities.scala 21:24]
  reg  _T_1795_1; // @[GameUtilities.scala 21:24]
  wire  _T_1797 = _T_1794_0 & _T_1795_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1800 = _T_1797 & _T_519; // @[SpriteBlender.scala 63:35]
  wire  _T_1801 = 7'h40 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_64 = _T_1800 & _T_1801; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_64 = io_datareader_64[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1806_0; // @[GameUtilities.scala 21:24]
  reg  _T_1806_1; // @[GameUtilities.scala 21:24]
  reg  _T_1807_0; // @[GameUtilities.scala 21:24]
  reg  _T_1807_1; // @[GameUtilities.scala 21:24]
  wire  _T_1809 = _T_1806_0 & _T_1807_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1812 = _T_1809 & _T_527; // @[SpriteBlender.scala 63:35]
  wire  _T_1813 = 7'h41 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_65 = _T_1812 & _T_1813; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_65 = io_datareader_65[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1818_0; // @[GameUtilities.scala 21:24]
  reg  _T_1818_1; // @[GameUtilities.scala 21:24]
  reg  _T_1819_0; // @[GameUtilities.scala 21:24]
  reg  _T_1819_1; // @[GameUtilities.scala 21:24]
  wire  _T_1821 = _T_1818_0 & _T_1819_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1824 = _T_1821 & _T_535; // @[SpriteBlender.scala 63:35]
  wire  _T_1825 = 7'h42 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_66 = _T_1824 & _T_1825; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_66 = io_datareader_66[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1831_0; // @[GameUtilities.scala 21:24]
  reg  _T_1831_1; // @[GameUtilities.scala 21:24]
  wire  _T_1836 = _T_1831_0 & _T_543; // @[SpriteBlender.scala 63:35]
  wire  _T_1837 = 7'h43 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_67 = _T_1836 & _T_1837; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_67 = io_datareader_67[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1843_0; // @[GameUtilities.scala 21:24]
  reg  _T_1843_1; // @[GameUtilities.scala 21:24]
  wire  _T_1848 = _T_1843_0 & _T_551; // @[SpriteBlender.scala 63:35]
  wire  _T_1849 = 7'h44 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_68 = _T_1848 & _T_1849; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_68 = io_datareader_68[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1855_0; // @[GameUtilities.scala 21:24]
  reg  _T_1855_1; // @[GameUtilities.scala 21:24]
  wire  _T_1860 = _T_1855_0 & _T_559; // @[SpriteBlender.scala 63:35]
  wire  _T_1861 = 7'h45 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_69 = _T_1860 & _T_1861; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_69 = io_datareader_69[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1866_0; // @[GameUtilities.scala 21:24]
  reg  _T_1866_1; // @[GameUtilities.scala 21:24]
  reg  _T_1867_0; // @[GameUtilities.scala 21:24]
  reg  _T_1867_1; // @[GameUtilities.scala 21:24]
  wire  _T_1869 = _T_1866_0 & _T_1867_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1872 = _T_1869 & _T_567; // @[SpriteBlender.scala 63:35]
  wire  _T_1873 = 7'h46 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_70 = _T_1872 & _T_1873; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_70 = io_datareader_70[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1878_0; // @[GameUtilities.scala 21:24]
  reg  _T_1878_1; // @[GameUtilities.scala 21:24]
  reg  _T_1879_0; // @[GameUtilities.scala 21:24]
  reg  _T_1879_1; // @[GameUtilities.scala 21:24]
  wire  _T_1881 = _T_1878_0 & _T_1879_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1884 = _T_1881 & _T_575; // @[SpriteBlender.scala 63:35]
  wire  _T_1885 = 7'h47 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_71 = _T_1884 & _T_1885; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_71 = io_datareader_71[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1890_0; // @[GameUtilities.scala 21:24]
  reg  _T_1890_1; // @[GameUtilities.scala 21:24]
  reg  _T_1891_0; // @[GameUtilities.scala 21:24]
  reg  _T_1891_1; // @[GameUtilities.scala 21:24]
  wire  _T_1893 = _T_1890_0 & _T_1891_0; // @[SpriteBlender.scala 63:25]
  wire  _T_1896 = _T_1893 & _T_583; // @[SpriteBlender.scala 63:35]
  wire  _T_1897 = 7'h48 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_72 = _T_1896 & _T_1897; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_72 = io_datareader_72[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1903_0; // @[GameUtilities.scala 21:24]
  reg  _T_1903_1; // @[GameUtilities.scala 21:24]
  wire  _T_1908 = _T_1903_0 & _T_591; // @[SpriteBlender.scala 63:35]
  wire  _T_1909 = 7'h49 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_73 = _T_1908 & _T_1909; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_73 = io_datareader_73[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1915_0; // @[GameUtilities.scala 21:24]
  reg  _T_1915_1; // @[GameUtilities.scala 21:24]
  wire  _T_1920 = _T_1915_0 & _T_599; // @[SpriteBlender.scala 63:35]
  wire  _T_1921 = 7'h4a != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_74 = _T_1920 & _T_1921; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_74 = io_datareader_74[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1927_0; // @[GameUtilities.scala 21:24]
  reg  _T_1927_1; // @[GameUtilities.scala 21:24]
  wire  _T_1932 = _T_1927_0 & _T_607; // @[SpriteBlender.scala 63:35]
  wire  _T_1933 = 7'h4b != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_75 = _T_1932 & _T_1933; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_75 = io_datareader_75[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1939_0; // @[GameUtilities.scala 21:24]
  reg  _T_1939_1; // @[GameUtilities.scala 21:24]
  wire  _T_1944 = _T_1939_0 & _T_615; // @[SpriteBlender.scala 63:35]
  wire  _T_1945 = 7'h4c != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_76 = _T_1944 & _T_1945; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_76 = io_datareader_76[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1951_0; // @[GameUtilities.scala 21:24]
  reg  _T_1951_1; // @[GameUtilities.scala 21:24]
  wire  _T_1956 = _T_1951_0 & _T_623; // @[SpriteBlender.scala 63:35]
  wire  _T_1957 = 7'h4d != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_77 = _T_1956 & _T_1957; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_77 = io_datareader_77[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1963_0; // @[GameUtilities.scala 21:24]
  reg  _T_1963_1; // @[GameUtilities.scala 21:24]
  wire  _T_1968 = _T_1963_0 & _T_631; // @[SpriteBlender.scala 63:35]
  wire  _T_1969 = 7'h4e != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_78 = _T_1968 & _T_1969; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_78 = io_datareader_78[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1975_0; // @[GameUtilities.scala 21:24]
  reg  _T_1975_1; // @[GameUtilities.scala 21:24]
  wire  _T_1980 = _T_1975_0 & _T_639; // @[SpriteBlender.scala 63:35]
  wire  _T_1981 = 7'h4f != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_79 = _T_1980 & _T_1981; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_79 = io_datareader_79[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1987_0; // @[GameUtilities.scala 21:24]
  reg  _T_1987_1; // @[GameUtilities.scala 21:24]
  wire  _T_1992 = _T_1987_0 & _T_647; // @[SpriteBlender.scala 63:35]
  wire  _T_1993 = 7'h50 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_80 = _T_1992 & _T_1993; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_80 = io_datareader_80[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_1999_0; // @[GameUtilities.scala 21:24]
  reg  _T_1999_1; // @[GameUtilities.scala 21:24]
  wire  _T_2004 = _T_1999_0 & _T_655; // @[SpriteBlender.scala 63:35]
  wire  _T_2005 = 7'h51 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_81 = _T_2004 & _T_2005; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_81 = io_datareader_81[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2011_0; // @[GameUtilities.scala 21:24]
  reg  _T_2011_1; // @[GameUtilities.scala 21:24]
  wire  _T_2016 = _T_2011_0 & _T_663; // @[SpriteBlender.scala 63:35]
  wire  _T_2017 = 7'h52 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_82 = _T_2016 & _T_2017; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_82 = io_datareader_82[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2023_0; // @[GameUtilities.scala 21:24]
  reg  _T_2023_1; // @[GameUtilities.scala 21:24]
  wire  _T_2028 = _T_2023_0 & _T_671; // @[SpriteBlender.scala 63:35]
  wire  _T_2029 = 7'h53 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_83 = _T_2028 & _T_2029; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_83 = io_datareader_83[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2035_0; // @[GameUtilities.scala 21:24]
  reg  _T_2035_1; // @[GameUtilities.scala 21:24]
  wire  _T_2040 = _T_2035_0 & _T_679; // @[SpriteBlender.scala 63:35]
  wire  _T_2041 = 7'h54 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_84 = _T_2040 & _T_2041; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_84 = io_datareader_84[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2047_0; // @[GameUtilities.scala 21:24]
  reg  _T_2047_1; // @[GameUtilities.scala 21:24]
  wire  _T_2052 = _T_2047_0 & _T_687; // @[SpriteBlender.scala 63:35]
  wire  _T_2053 = 7'h55 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_85 = _T_2052 & _T_2053; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_85 = io_datareader_85[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2059_0; // @[GameUtilities.scala 21:24]
  reg  _T_2059_1; // @[GameUtilities.scala 21:24]
  wire  _T_2064 = _T_2059_0 & _T_695; // @[SpriteBlender.scala 63:35]
  wire  _T_2065 = 7'h56 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_86 = _T_2064 & _T_2065; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_86 = io_datareader_86[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2071_0; // @[GameUtilities.scala 21:24]
  reg  _T_2071_1; // @[GameUtilities.scala 21:24]
  wire  _T_2076 = _T_2071_0 & _T_703; // @[SpriteBlender.scala 63:35]
  wire  _T_2077 = 7'h57 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_87 = _T_2076 & _T_2077; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_87 = io_datareader_87[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2083_0; // @[GameUtilities.scala 21:24]
  reg  _T_2083_1; // @[GameUtilities.scala 21:24]
  wire  _T_2088 = _T_2083_0 & _T_711; // @[SpriteBlender.scala 63:35]
  wire  _T_2089 = 7'h58 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_88 = _T_2088 & _T_2089; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_88 = io_datareader_88[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2095_0; // @[GameUtilities.scala 21:24]
  reg  _T_2095_1; // @[GameUtilities.scala 21:24]
  wire  _T_2100 = _T_2095_0 & _T_719; // @[SpriteBlender.scala 63:35]
  wire  _T_2101 = 7'h59 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_89 = _T_2100 & _T_2101; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_89 = io_datareader_89[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2107_0; // @[GameUtilities.scala 21:24]
  reg  _T_2107_1; // @[GameUtilities.scala 21:24]
  wire  _T_2112 = _T_2107_0 & _T_727; // @[SpriteBlender.scala 63:35]
  wire  _T_2113 = 7'h5a != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_90 = _T_2112 & _T_2113; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_90 = io_datareader_90[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2119_0; // @[GameUtilities.scala 21:24]
  reg  _T_2119_1; // @[GameUtilities.scala 21:24]
  wire  _T_2124 = _T_2119_0 & _T_735; // @[SpriteBlender.scala 63:35]
  wire  _T_2125 = 7'h5b != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_91 = _T_2124 & _T_2125; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_91 = io_datareader_91[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2131_0; // @[GameUtilities.scala 21:24]
  reg  _T_2131_1; // @[GameUtilities.scala 21:24]
  wire  _T_2136 = _T_2131_0 & _T_743; // @[SpriteBlender.scala 63:35]
  wire  _T_2137 = 7'h5c != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_92 = _T_2136 & _T_2137; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_92 = io_datareader_92[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2143_0; // @[GameUtilities.scala 21:24]
  reg  _T_2143_1; // @[GameUtilities.scala 21:24]
  wire  _T_2148 = _T_2143_0 & _T_751; // @[SpriteBlender.scala 63:35]
  wire  _T_2149 = 7'h5d != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_93 = _T_2148 & _T_2149; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_93 = io_datareader_93[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2155_0; // @[GameUtilities.scala 21:24]
  reg  _T_2155_1; // @[GameUtilities.scala 21:24]
  wire  _T_2160 = _T_2155_0 & _T_759; // @[SpriteBlender.scala 63:35]
  wire  _T_2161 = 7'h5e != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_94 = _T_2160 & _T_2161; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_94 = io_datareader_94[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2167_0; // @[GameUtilities.scala 21:24]
  reg  _T_2167_1; // @[GameUtilities.scala 21:24]
  wire  _T_2172 = _T_2167_0 & _T_767; // @[SpriteBlender.scala 63:35]
  wire  _T_2173 = 7'h5f != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_95 = _T_2172 & _T_2173; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_95 = io_datareader_95[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2179_0; // @[GameUtilities.scala 21:24]
  reg  _T_2179_1; // @[GameUtilities.scala 21:24]
  wire  _T_2184 = _T_2179_0 & _T_775; // @[SpriteBlender.scala 63:35]
  wire  _T_2185 = 7'h60 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_96 = _T_2184 & _T_2185; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_96 = io_datareader_96[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2191_0; // @[GameUtilities.scala 21:24]
  reg  _T_2191_1; // @[GameUtilities.scala 21:24]
  wire  _T_2196 = _T_2191_0 & _T_783; // @[SpriteBlender.scala 63:35]
  wire  _T_2197 = 7'h61 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_97 = _T_2196 & _T_2197; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_97 = io_datareader_97[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2203_0; // @[GameUtilities.scala 21:24]
  reg  _T_2203_1; // @[GameUtilities.scala 21:24]
  wire  _T_2208 = _T_2203_0 & _T_791; // @[SpriteBlender.scala 63:35]
  wire  _T_2209 = 7'h62 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_98 = _T_2208 & _T_2209; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_98 = io_datareader_98[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2215_0; // @[GameUtilities.scala 21:24]
  reg  _T_2215_1; // @[GameUtilities.scala 21:24]
  wire  _T_2220 = _T_2215_0 & _T_799; // @[SpriteBlender.scala 63:35]
  wire  _T_2221 = 7'h63 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_99 = _T_2220 & _T_2221; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_99 = io_datareader_99[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2227_0; // @[GameUtilities.scala 21:24]
  reg  _T_2227_1; // @[GameUtilities.scala 21:24]
  wire  _T_2232 = _T_2227_0 & _T_807; // @[SpriteBlender.scala 63:35]
  wire  _T_2233 = 7'h64 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_100 = _T_2232 & _T_2233; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_100 = io_datareader_100[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2239_0; // @[GameUtilities.scala 21:24]
  reg  _T_2239_1; // @[GameUtilities.scala 21:24]
  wire  _T_2244 = _T_2239_0 & _T_815; // @[SpriteBlender.scala 63:35]
  wire  _T_2245 = 7'h65 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_101 = _T_2244 & _T_2245; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_101 = io_datareader_101[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2251_0; // @[GameUtilities.scala 21:24]
  reg  _T_2251_1; // @[GameUtilities.scala 21:24]
  wire  _T_2256 = _T_2251_0 & _T_823; // @[SpriteBlender.scala 63:35]
  wire  _T_2257 = 7'h66 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_102 = _T_2256 & _T_2257; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_102 = io_datareader_102[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2263_0; // @[GameUtilities.scala 21:24]
  reg  _T_2263_1; // @[GameUtilities.scala 21:24]
  wire  _T_2268 = _T_2263_0 & _T_831; // @[SpriteBlender.scala 63:35]
  wire  _T_2269 = 7'h67 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_103 = _T_2268 & _T_2269; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_103 = io_datareader_103[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2275_0; // @[GameUtilities.scala 21:24]
  reg  _T_2275_1; // @[GameUtilities.scala 21:24]
  wire  _T_2280 = _T_2275_0 & _T_839; // @[SpriteBlender.scala 63:35]
  wire  _T_2281 = 7'h68 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_104 = _T_2280 & _T_2281; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_104 = io_datareader_104[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2287_0; // @[GameUtilities.scala 21:24]
  reg  _T_2287_1; // @[GameUtilities.scala 21:24]
  wire  _T_2292 = _T_2287_0 & _T_847; // @[SpriteBlender.scala 63:35]
  wire  _T_2293 = 7'h69 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_105 = _T_2292 & _T_2293; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_105 = io_datareader_105[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2299_0; // @[GameUtilities.scala 21:24]
  reg  _T_2299_1; // @[GameUtilities.scala 21:24]
  wire  _T_2304 = _T_2299_0 & _T_855; // @[SpriteBlender.scala 63:35]
  wire  _T_2305 = 7'h6a != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_106 = _T_2304 & _T_2305; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_106 = io_datareader_106[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2311_0; // @[GameUtilities.scala 21:24]
  reg  _T_2311_1; // @[GameUtilities.scala 21:24]
  wire  _T_2316 = _T_2311_0 & _T_863; // @[SpriteBlender.scala 63:35]
  wire  _T_2317 = 7'h6b != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_107 = _T_2316 & _T_2317; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_107 = io_datareader_107[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2323_0; // @[GameUtilities.scala 21:24]
  reg  _T_2323_1; // @[GameUtilities.scala 21:24]
  wire  _T_2328 = _T_2323_0 & _T_871; // @[SpriteBlender.scala 63:35]
  wire  _T_2329 = 7'h6c != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_108 = _T_2328 & _T_2329; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_108 = io_datareader_108[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2335_0; // @[GameUtilities.scala 21:24]
  reg  _T_2335_1; // @[GameUtilities.scala 21:24]
  wire  _T_2340 = _T_2335_0 & _T_879; // @[SpriteBlender.scala 63:35]
  wire  _T_2341 = 7'h6d != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_109 = _T_2340 & _T_2341; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_109 = io_datareader_109[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2347_0; // @[GameUtilities.scala 21:24]
  reg  _T_2347_1; // @[GameUtilities.scala 21:24]
  wire  _T_2352 = _T_2347_0 & _T_887; // @[SpriteBlender.scala 63:35]
  wire  _T_2353 = 7'h6e != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_110 = _T_2352 & _T_2353; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_110 = io_datareader_110[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2359_0; // @[GameUtilities.scala 21:24]
  reg  _T_2359_1; // @[GameUtilities.scala 21:24]
  wire  _T_2364 = _T_2359_0 & _T_895; // @[SpriteBlender.scala 63:35]
  wire  _T_2365 = 7'h6f != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_111 = _T_2364 & _T_2365; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_111 = io_datareader_111[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2371_0; // @[GameUtilities.scala 21:24]
  reg  _T_2371_1; // @[GameUtilities.scala 21:24]
  wire  _T_2376 = _T_2371_0 & _T_903; // @[SpriteBlender.scala 63:35]
  wire  _T_2377 = 7'h70 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_112 = _T_2376 & _T_2377; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_112 = io_datareader_112[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2383_0; // @[GameUtilities.scala 21:24]
  reg  _T_2383_1; // @[GameUtilities.scala 21:24]
  wire  _T_2388 = _T_2383_0 & _T_911; // @[SpriteBlender.scala 63:35]
  wire  _T_2389 = 7'h71 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_113 = _T_2388 & _T_2389; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_113 = io_datareader_113[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2395_0; // @[GameUtilities.scala 21:24]
  reg  _T_2395_1; // @[GameUtilities.scala 21:24]
  wire  _T_2400 = _T_2395_0 & _T_919; // @[SpriteBlender.scala 63:35]
  wire  _T_2401 = 7'h72 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_114 = _T_2400 & _T_2401; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_114 = io_datareader_114[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2407_0; // @[GameUtilities.scala 21:24]
  reg  _T_2407_1; // @[GameUtilities.scala 21:24]
  wire  _T_2412 = _T_2407_0 & _T_927; // @[SpriteBlender.scala 63:35]
  wire  _T_2413 = 7'h73 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_115 = _T_2412 & _T_2413; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_115 = io_datareader_115[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2419_0; // @[GameUtilities.scala 21:24]
  reg  _T_2419_1; // @[GameUtilities.scala 21:24]
  wire  _T_2424 = _T_2419_0 & _T_935; // @[SpriteBlender.scala 63:35]
  wire  _T_2425 = 7'h74 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_116 = _T_2424 & _T_2425; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_116 = io_datareader_116[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2431_0; // @[GameUtilities.scala 21:24]
  reg  _T_2431_1; // @[GameUtilities.scala 21:24]
  wire  _T_2436 = _T_2431_0 & _T_943; // @[SpriteBlender.scala 63:35]
  wire  _T_2437 = 7'h75 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_117 = _T_2436 & _T_2437; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_117 = io_datareader_117[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2443_0; // @[GameUtilities.scala 21:24]
  reg  _T_2443_1; // @[GameUtilities.scala 21:24]
  wire  _T_2448 = _T_2443_0 & _T_951; // @[SpriteBlender.scala 63:35]
  wire  _T_2449 = 7'h76 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_118 = _T_2448 & _T_2449; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_118 = io_datareader_118[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2455_0; // @[GameUtilities.scala 21:24]
  reg  _T_2455_1; // @[GameUtilities.scala 21:24]
  wire  _T_2460 = _T_2455_0 & _T_959; // @[SpriteBlender.scala 63:35]
  wire  _T_2461 = 7'h77 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_119 = _T_2460 & _T_2461; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_119 = io_datareader_119[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2467_0; // @[GameUtilities.scala 21:24]
  reg  _T_2467_1; // @[GameUtilities.scala 21:24]
  wire  _T_2472 = _T_2467_0 & _T_967; // @[SpriteBlender.scala 63:35]
  wire  _T_2473 = 7'h78 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_120 = _T_2472 & _T_2473; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_120 = io_datareader_120[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2479_0; // @[GameUtilities.scala 21:24]
  reg  _T_2479_1; // @[GameUtilities.scala 21:24]
  wire  _T_2484 = _T_2479_0 & _T_975; // @[SpriteBlender.scala 63:35]
  wire  _T_2485 = 7'h79 != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_121 = _T_2484 & _T_2485; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_121 = io_datareader_121[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2491_0; // @[GameUtilities.scala 21:24]
  reg  _T_2491_1; // @[GameUtilities.scala 21:24]
  wire  _T_2496 = _T_2491_0 & _T_983; // @[SpriteBlender.scala 63:35]
  wire  _T_2497 = 7'h7a != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_122 = _T_2496 & _T_2497; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_122 = io_datareader_122[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2503_0; // @[GameUtilities.scala 21:24]
  reg  _T_2503_1; // @[GameUtilities.scala 21:24]
  wire  _T_2508 = _T_2503_0 & _T_991; // @[SpriteBlender.scala 63:35]
  wire  _T_2509 = 7'h7b != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_123 = _T_2508 & _T_2509; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_123 = io_datareader_123[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2515_0; // @[GameUtilities.scala 21:24]
  reg  _T_2515_1; // @[GameUtilities.scala 21:24]
  wire  _T_2520 = _T_2515_0 & _T_999; // @[SpriteBlender.scala 63:35]
  wire  _T_2521 = 7'h7c != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_124 = _T_2520 & _T_2521; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_124 = io_datareader_124[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2527_0; // @[GameUtilities.scala 21:24]
  reg  _T_2527_1; // @[GameUtilities.scala 21:24]
  wire  _T_2532 = _T_2527_0 & _T_1007; // @[SpriteBlender.scala 63:35]
  wire  _T_2533 = 7'h7d != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_125 = _T_2532 & _T_2533; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_125 = io_datareader_125[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2539_0; // @[GameUtilities.scala 21:24]
  reg  _T_2539_1; // @[GameUtilities.scala 21:24]
  wire  _T_2544 = _T_2539_0 & _T_1015; // @[SpriteBlender.scala 63:35]
  wire  _T_2545 = 7'h7e != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_126 = _T_2544 & _T_2545; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_126 = io_datareader_126[5:0]; // @[SpriteBlender.scala 65:44]
  reg  _T_2551_0; // @[GameUtilities.scala 21:24]
  reg  _T_2551_1; // @[GameUtilities.scala 21:24]
  wire  _T_2556 = _T_2551_0 & _T_1023; // @[SpriteBlender.scala 63:35]
  wire  _T_2557 = 7'h7f != multiHotPriortyReductionTree_io_indexOutput; // @[SpriteBlender.scala 63:63]
  wire  secondSpriteValids_127 = _T_2556 & _T_2557; // @[SpriteBlender.scala 63:55]
  wire [5:0] secondSpriteCandidates_127 = io_datareader_127[5:0]; // @[SpriteBlender.scala 65:44]
  wire [5:0] _T_2562 = secondSpriteValids_126 ? secondSpriteCandidates_126 : secondSpriteCandidates_127; // @[Mux.scala 47:69]
  wire [5:0] _T_2563 = secondSpriteValids_125 ? secondSpriteCandidates_125 : _T_2562; // @[Mux.scala 47:69]
  wire [5:0] _T_2564 = secondSpriteValids_124 ? secondSpriteCandidates_124 : _T_2563; // @[Mux.scala 47:69]
  wire [5:0] _T_2565 = secondSpriteValids_123 ? secondSpriteCandidates_123 : _T_2564; // @[Mux.scala 47:69]
  wire [5:0] _T_2566 = secondSpriteValids_122 ? secondSpriteCandidates_122 : _T_2565; // @[Mux.scala 47:69]
  wire [5:0] _T_2567 = secondSpriteValids_121 ? secondSpriteCandidates_121 : _T_2566; // @[Mux.scala 47:69]
  wire [5:0] _T_2568 = secondSpriteValids_120 ? secondSpriteCandidates_120 : _T_2567; // @[Mux.scala 47:69]
  wire [5:0] _T_2569 = secondSpriteValids_119 ? secondSpriteCandidates_119 : _T_2568; // @[Mux.scala 47:69]
  wire [5:0] _T_2570 = secondSpriteValids_118 ? secondSpriteCandidates_118 : _T_2569; // @[Mux.scala 47:69]
  wire [5:0] _T_2571 = secondSpriteValids_117 ? secondSpriteCandidates_117 : _T_2570; // @[Mux.scala 47:69]
  wire [5:0] _T_2572 = secondSpriteValids_116 ? secondSpriteCandidates_116 : _T_2571; // @[Mux.scala 47:69]
  wire [5:0] _T_2573 = secondSpriteValids_115 ? secondSpriteCandidates_115 : _T_2572; // @[Mux.scala 47:69]
  wire [5:0] _T_2574 = secondSpriteValids_114 ? secondSpriteCandidates_114 : _T_2573; // @[Mux.scala 47:69]
  wire [5:0] _T_2575 = secondSpriteValids_113 ? secondSpriteCandidates_113 : _T_2574; // @[Mux.scala 47:69]
  wire [5:0] _T_2576 = secondSpriteValids_112 ? secondSpriteCandidates_112 : _T_2575; // @[Mux.scala 47:69]
  wire [5:0] _T_2577 = secondSpriteValids_111 ? secondSpriteCandidates_111 : _T_2576; // @[Mux.scala 47:69]
  wire [5:0] _T_2578 = secondSpriteValids_110 ? secondSpriteCandidates_110 : _T_2577; // @[Mux.scala 47:69]
  wire [5:0] _T_2579 = secondSpriteValids_109 ? secondSpriteCandidates_109 : _T_2578; // @[Mux.scala 47:69]
  wire [5:0] _T_2580 = secondSpriteValids_108 ? secondSpriteCandidates_108 : _T_2579; // @[Mux.scala 47:69]
  wire [5:0] _T_2581 = secondSpriteValids_107 ? secondSpriteCandidates_107 : _T_2580; // @[Mux.scala 47:69]
  wire [5:0] _T_2582 = secondSpriteValids_106 ? secondSpriteCandidates_106 : _T_2581; // @[Mux.scala 47:69]
  wire [5:0] _T_2583 = secondSpriteValids_105 ? secondSpriteCandidates_105 : _T_2582; // @[Mux.scala 47:69]
  wire [5:0] _T_2584 = secondSpriteValids_104 ? secondSpriteCandidates_104 : _T_2583; // @[Mux.scala 47:69]
  wire [5:0] _T_2585 = secondSpriteValids_103 ? secondSpriteCandidates_103 : _T_2584; // @[Mux.scala 47:69]
  wire [5:0] _T_2586 = secondSpriteValids_102 ? secondSpriteCandidates_102 : _T_2585; // @[Mux.scala 47:69]
  wire [5:0] _T_2587 = secondSpriteValids_101 ? secondSpriteCandidates_101 : _T_2586; // @[Mux.scala 47:69]
  wire [5:0] _T_2588 = secondSpriteValids_100 ? secondSpriteCandidates_100 : _T_2587; // @[Mux.scala 47:69]
  wire [5:0] _T_2589 = secondSpriteValids_99 ? secondSpriteCandidates_99 : _T_2588; // @[Mux.scala 47:69]
  wire [5:0] _T_2590 = secondSpriteValids_98 ? secondSpriteCandidates_98 : _T_2589; // @[Mux.scala 47:69]
  wire [5:0] _T_2591 = secondSpriteValids_97 ? secondSpriteCandidates_97 : _T_2590; // @[Mux.scala 47:69]
  wire [5:0] _T_2592 = secondSpriteValids_96 ? secondSpriteCandidates_96 : _T_2591; // @[Mux.scala 47:69]
  wire [5:0] _T_2593 = secondSpriteValids_95 ? secondSpriteCandidates_95 : _T_2592; // @[Mux.scala 47:69]
  wire [5:0] _T_2594 = secondSpriteValids_94 ? secondSpriteCandidates_94 : _T_2593; // @[Mux.scala 47:69]
  wire [5:0] _T_2595 = secondSpriteValids_93 ? secondSpriteCandidates_93 : _T_2594; // @[Mux.scala 47:69]
  wire [5:0] _T_2596 = secondSpriteValids_92 ? secondSpriteCandidates_92 : _T_2595; // @[Mux.scala 47:69]
  wire [5:0] _T_2597 = secondSpriteValids_91 ? secondSpriteCandidates_91 : _T_2596; // @[Mux.scala 47:69]
  wire [5:0] _T_2598 = secondSpriteValids_90 ? secondSpriteCandidates_90 : _T_2597; // @[Mux.scala 47:69]
  wire [5:0] _T_2599 = secondSpriteValids_89 ? secondSpriteCandidates_89 : _T_2598; // @[Mux.scala 47:69]
  wire [5:0] _T_2600 = secondSpriteValids_88 ? secondSpriteCandidates_88 : _T_2599; // @[Mux.scala 47:69]
  wire [5:0] _T_2601 = secondSpriteValids_87 ? secondSpriteCandidates_87 : _T_2600; // @[Mux.scala 47:69]
  wire [5:0] _T_2602 = secondSpriteValids_86 ? secondSpriteCandidates_86 : _T_2601; // @[Mux.scala 47:69]
  wire [5:0] _T_2603 = secondSpriteValids_85 ? secondSpriteCandidates_85 : _T_2602; // @[Mux.scala 47:69]
  wire [5:0] _T_2604 = secondSpriteValids_84 ? secondSpriteCandidates_84 : _T_2603; // @[Mux.scala 47:69]
  wire [5:0] _T_2605 = secondSpriteValids_83 ? secondSpriteCandidates_83 : _T_2604; // @[Mux.scala 47:69]
  wire [5:0] _T_2606 = secondSpriteValids_82 ? secondSpriteCandidates_82 : _T_2605; // @[Mux.scala 47:69]
  wire [5:0] _T_2607 = secondSpriteValids_81 ? secondSpriteCandidates_81 : _T_2606; // @[Mux.scala 47:69]
  wire [5:0] _T_2608 = secondSpriteValids_80 ? secondSpriteCandidates_80 : _T_2607; // @[Mux.scala 47:69]
  wire [5:0] _T_2609 = secondSpriteValids_79 ? secondSpriteCandidates_79 : _T_2608; // @[Mux.scala 47:69]
  wire [5:0] _T_2610 = secondSpriteValids_78 ? secondSpriteCandidates_78 : _T_2609; // @[Mux.scala 47:69]
  wire [5:0] _T_2611 = secondSpriteValids_77 ? secondSpriteCandidates_77 : _T_2610; // @[Mux.scala 47:69]
  wire [5:0] _T_2612 = secondSpriteValids_76 ? secondSpriteCandidates_76 : _T_2611; // @[Mux.scala 47:69]
  wire [5:0] _T_2613 = secondSpriteValids_75 ? secondSpriteCandidates_75 : _T_2612; // @[Mux.scala 47:69]
  wire [5:0] _T_2614 = secondSpriteValids_74 ? secondSpriteCandidates_74 : _T_2613; // @[Mux.scala 47:69]
  wire [5:0] _T_2615 = secondSpriteValids_73 ? secondSpriteCandidates_73 : _T_2614; // @[Mux.scala 47:69]
  wire [5:0] _T_2616 = secondSpriteValids_72 ? secondSpriteCandidates_72 : _T_2615; // @[Mux.scala 47:69]
  wire [5:0] _T_2617 = secondSpriteValids_71 ? secondSpriteCandidates_71 : _T_2616; // @[Mux.scala 47:69]
  wire [5:0] _T_2618 = secondSpriteValids_70 ? secondSpriteCandidates_70 : _T_2617; // @[Mux.scala 47:69]
  wire [5:0] _T_2619 = secondSpriteValids_69 ? secondSpriteCandidates_69 : _T_2618; // @[Mux.scala 47:69]
  wire [5:0] _T_2620 = secondSpriteValids_68 ? secondSpriteCandidates_68 : _T_2619; // @[Mux.scala 47:69]
  wire [5:0] _T_2621 = secondSpriteValids_67 ? secondSpriteCandidates_67 : _T_2620; // @[Mux.scala 47:69]
  wire [5:0] _T_2622 = secondSpriteValids_66 ? secondSpriteCandidates_66 : _T_2621; // @[Mux.scala 47:69]
  wire [5:0] _T_2623 = secondSpriteValids_65 ? secondSpriteCandidates_65 : _T_2622; // @[Mux.scala 47:69]
  wire [5:0] _T_2624 = secondSpriteValids_64 ? secondSpriteCandidates_64 : _T_2623; // @[Mux.scala 47:69]
  wire [5:0] _T_2625 = secondSpriteValids_63 ? secondSpriteCandidates_63 : _T_2624; // @[Mux.scala 47:69]
  wire [5:0] _T_2626 = secondSpriteValids_62 ? secondSpriteCandidates_62 : _T_2625; // @[Mux.scala 47:69]
  wire [5:0] _T_2627 = secondSpriteValids_61 ? secondSpriteCandidates_61 : _T_2626; // @[Mux.scala 47:69]
  wire [5:0] _T_2628 = secondSpriteValids_60 ? secondSpriteCandidates_60 : _T_2627; // @[Mux.scala 47:69]
  wire [5:0] _T_2629 = secondSpriteValids_59 ? secondSpriteCandidates_59 : _T_2628; // @[Mux.scala 47:69]
  wire [5:0] _T_2630 = secondSpriteValids_58 ? secondSpriteCandidates_58 : _T_2629; // @[Mux.scala 47:69]
  wire [5:0] _T_2631 = secondSpriteValids_57 ? secondSpriteCandidates_57 : _T_2630; // @[Mux.scala 47:69]
  wire [5:0] _T_2632 = secondSpriteValids_56 ? secondSpriteCandidates_56 : _T_2631; // @[Mux.scala 47:69]
  wire [5:0] _T_2633 = secondSpriteValids_55 ? secondSpriteCandidates_55 : _T_2632; // @[Mux.scala 47:69]
  wire [5:0] _T_2634 = secondSpriteValids_54 ? secondSpriteCandidates_54 : _T_2633; // @[Mux.scala 47:69]
  wire [5:0] _T_2635 = secondSpriteValids_53 ? secondSpriteCandidates_53 : _T_2634; // @[Mux.scala 47:69]
  wire [5:0] _T_2636 = secondSpriteValids_52 ? secondSpriteCandidates_52 : _T_2635; // @[Mux.scala 47:69]
  wire [5:0] _T_2637 = secondSpriteValids_51 ? secondSpriteCandidates_51 : _T_2636; // @[Mux.scala 47:69]
  wire [5:0] _T_2638 = secondSpriteValids_50 ? secondSpriteCandidates_50 : _T_2637; // @[Mux.scala 47:69]
  wire [5:0] _T_2639 = secondSpriteValids_49 ? secondSpriteCandidates_49 : _T_2638; // @[Mux.scala 47:69]
  wire [5:0] _T_2640 = secondSpriteValids_48 ? secondSpriteCandidates_48 : _T_2639; // @[Mux.scala 47:69]
  wire [5:0] _T_2641 = secondSpriteValids_47 ? secondSpriteCandidates_47 : _T_2640; // @[Mux.scala 47:69]
  wire [5:0] _T_2642 = secondSpriteValids_46 ? secondSpriteCandidates_46 : _T_2641; // @[Mux.scala 47:69]
  wire [5:0] _T_2643 = secondSpriteValids_45 ? secondSpriteCandidates_45 : _T_2642; // @[Mux.scala 47:69]
  wire [5:0] _T_2644 = secondSpriteValids_44 ? secondSpriteCandidates_44 : _T_2643; // @[Mux.scala 47:69]
  wire [5:0] _T_2645 = secondSpriteValids_43 ? secondSpriteCandidates_43 : _T_2644; // @[Mux.scala 47:69]
  wire [5:0] _T_2646 = secondSpriteValids_42 ? secondSpriteCandidates_42 : _T_2645; // @[Mux.scala 47:69]
  wire [5:0] _T_2647 = secondSpriteValids_41 ? secondSpriteCandidates_41 : _T_2646; // @[Mux.scala 47:69]
  wire [5:0] _T_2648 = secondSpriteValids_40 ? secondSpriteCandidates_40 : _T_2647; // @[Mux.scala 47:69]
  wire [5:0] _T_2649 = secondSpriteValids_39 ? secondSpriteCandidates_39 : _T_2648; // @[Mux.scala 47:69]
  wire [5:0] _T_2650 = secondSpriteValids_38 ? secondSpriteCandidates_38 : _T_2649; // @[Mux.scala 47:69]
  wire [5:0] _T_2651 = secondSpriteValids_37 ? secondSpriteCandidates_37 : _T_2650; // @[Mux.scala 47:69]
  wire [5:0] _T_2652 = secondSpriteValids_36 ? secondSpriteCandidates_36 : _T_2651; // @[Mux.scala 47:69]
  wire [5:0] _T_2653 = secondSpriteValids_35 ? secondSpriteCandidates_35 : _T_2652; // @[Mux.scala 47:69]
  wire [5:0] _T_2654 = secondSpriteValids_34 ? secondSpriteCandidates_34 : _T_2653; // @[Mux.scala 47:69]
  wire [5:0] _T_2655 = secondSpriteValids_33 ? secondSpriteCandidates_33 : _T_2654; // @[Mux.scala 47:69]
  wire [5:0] _T_2656 = secondSpriteValids_32 ? secondSpriteCandidates_32 : _T_2655; // @[Mux.scala 47:69]
  wire [5:0] _T_2657 = secondSpriteValids_31 ? secondSpriteCandidates_31 : _T_2656; // @[Mux.scala 47:69]
  wire [5:0] _T_2658 = secondSpriteValids_30 ? secondSpriteCandidates_30 : _T_2657; // @[Mux.scala 47:69]
  wire [5:0] _T_2659 = secondSpriteValids_29 ? secondSpriteCandidates_29 : _T_2658; // @[Mux.scala 47:69]
  wire [5:0] _T_2660 = secondSpriteValids_28 ? secondSpriteCandidates_28 : _T_2659; // @[Mux.scala 47:69]
  wire [5:0] _T_2661 = secondSpriteValids_27 ? secondSpriteCandidates_27 : _T_2660; // @[Mux.scala 47:69]
  wire [5:0] _T_2662 = secondSpriteValids_26 ? secondSpriteCandidates_26 : _T_2661; // @[Mux.scala 47:69]
  wire [5:0] _T_2663 = secondSpriteValids_25 ? secondSpriteCandidates_25 : _T_2662; // @[Mux.scala 47:69]
  wire [5:0] _T_2664 = secondSpriteValids_24 ? secondSpriteCandidates_24 : _T_2663; // @[Mux.scala 47:69]
  wire [5:0] _T_2665 = secondSpriteValids_23 ? secondSpriteCandidates_23 : _T_2664; // @[Mux.scala 47:69]
  wire [5:0] _T_2666 = secondSpriteValids_22 ? secondSpriteCandidates_22 : _T_2665; // @[Mux.scala 47:69]
  wire [5:0] _T_2667 = secondSpriteValids_21 ? secondSpriteCandidates_21 : _T_2666; // @[Mux.scala 47:69]
  wire [5:0] _T_2668 = secondSpriteValids_20 ? secondSpriteCandidates_20 : _T_2667; // @[Mux.scala 47:69]
  wire [5:0] _T_2669 = secondSpriteValids_19 ? secondSpriteCandidates_19 : _T_2668; // @[Mux.scala 47:69]
  wire [5:0] _T_2670 = secondSpriteValids_18 ? secondSpriteCandidates_18 : _T_2669; // @[Mux.scala 47:69]
  wire [5:0] _T_2671 = secondSpriteValids_17 ? secondSpriteCandidates_17 : _T_2670; // @[Mux.scala 47:69]
  wire [5:0] _T_2672 = secondSpriteValids_16 ? secondSpriteCandidates_16 : _T_2671; // @[Mux.scala 47:69]
  wire [5:0] _T_2673 = secondSpriteValids_15 ? secondSpriteCandidates_15 : _T_2672; // @[Mux.scala 47:69]
  wire [5:0] _T_2674 = secondSpriteValids_14 ? secondSpriteCandidates_14 : _T_2673; // @[Mux.scala 47:69]
  wire [5:0] _T_2675 = secondSpriteValids_13 ? secondSpriteCandidates_13 : _T_2674; // @[Mux.scala 47:69]
  wire [5:0] _T_2676 = secondSpriteValids_12 ? secondSpriteCandidates_12 : _T_2675; // @[Mux.scala 47:69]
  wire [5:0] _T_2677 = secondSpriteValids_11 ? secondSpriteCandidates_11 : _T_2676; // @[Mux.scala 47:69]
  wire [5:0] _T_2678 = secondSpriteValids_10 ? secondSpriteCandidates_10 : _T_2677; // @[Mux.scala 47:69]
  wire [5:0] _T_2679 = secondSpriteValids_9 ? secondSpriteCandidates_9 : _T_2678; // @[Mux.scala 47:69]
  wire [5:0] _T_2680 = secondSpriteValids_8 ? secondSpriteCandidates_8 : _T_2679; // @[Mux.scala 47:69]
  wire [5:0] _T_2681 = secondSpriteValids_7 ? secondSpriteCandidates_7 : _T_2680; // @[Mux.scala 47:69]
  wire [5:0] _T_2682 = secondSpriteValids_6 ? secondSpriteCandidates_6 : _T_2681; // @[Mux.scala 47:69]
  wire [5:0] _T_2683 = secondSpriteValids_5 ? secondSpriteCandidates_5 : _T_2682; // @[Mux.scala 47:69]
  wire [5:0] _T_2684 = secondSpriteValids_4 ? secondSpriteCandidates_4 : _T_2683; // @[Mux.scala 47:69]
  wire [5:0] _T_2685 = secondSpriteValids_3 ? secondSpriteCandidates_3 : _T_2684; // @[Mux.scala 47:69]
  wire [5:0] _T_2686 = secondSpriteValids_2 ? secondSpriteCandidates_2 : _T_2685; // @[Mux.scala 47:69]
  wire [5:0] _T_2687 = secondSpriteValids_1 ? secondSpriteCandidates_1 : _T_2686; // @[Mux.scala 47:69]
  wire [5:0] secondTopSpriteColor = secondSpriteValids_0 ? secondSpriteCandidates_0 : _T_2687; // @[Mux.scala 47:69]
  wire  _T_2816 = secondSpriteValids_0 | secondSpriteValids_1; // @[SpriteBlender.scala 81:55]
  wire  _T_2817 = _T_2816 | secondSpriteValids_2; // @[SpriteBlender.scala 81:55]
  wire  _T_2818 = _T_2817 | secondSpriteValids_3; // @[SpriteBlender.scala 81:55]
  wire  _T_2819 = _T_2818 | secondSpriteValids_4; // @[SpriteBlender.scala 81:55]
  wire  _T_2820 = _T_2819 | secondSpriteValids_5; // @[SpriteBlender.scala 81:55]
  wire  _T_2821 = _T_2820 | secondSpriteValids_6; // @[SpriteBlender.scala 81:55]
  wire  _T_2822 = _T_2821 | secondSpriteValids_7; // @[SpriteBlender.scala 81:55]
  wire  _T_2823 = _T_2822 | secondSpriteValids_8; // @[SpriteBlender.scala 81:55]
  wire  _T_2824 = _T_2823 | secondSpriteValids_9; // @[SpriteBlender.scala 81:55]
  wire  _T_2825 = _T_2824 | secondSpriteValids_10; // @[SpriteBlender.scala 81:55]
  wire  _T_2826 = _T_2825 | secondSpriteValids_11; // @[SpriteBlender.scala 81:55]
  wire  _T_2827 = _T_2826 | secondSpriteValids_12; // @[SpriteBlender.scala 81:55]
  wire  _T_2828 = _T_2827 | secondSpriteValids_13; // @[SpriteBlender.scala 81:55]
  wire  _T_2829 = _T_2828 | secondSpriteValids_14; // @[SpriteBlender.scala 81:55]
  wire  _T_2830 = _T_2829 | secondSpriteValids_15; // @[SpriteBlender.scala 81:55]
  wire  _T_2831 = _T_2830 | secondSpriteValids_16; // @[SpriteBlender.scala 81:55]
  wire  _T_2832 = _T_2831 | secondSpriteValids_17; // @[SpriteBlender.scala 81:55]
  wire  _T_2833 = _T_2832 | secondSpriteValids_18; // @[SpriteBlender.scala 81:55]
  wire  _T_2834 = _T_2833 | secondSpriteValids_19; // @[SpriteBlender.scala 81:55]
  wire  _T_2835 = _T_2834 | secondSpriteValids_20; // @[SpriteBlender.scala 81:55]
  wire  _T_2836 = _T_2835 | secondSpriteValids_21; // @[SpriteBlender.scala 81:55]
  wire  _T_2837 = _T_2836 | secondSpriteValids_22; // @[SpriteBlender.scala 81:55]
  wire  _T_2838 = _T_2837 | secondSpriteValids_23; // @[SpriteBlender.scala 81:55]
  wire  _T_2839 = _T_2838 | secondSpriteValids_24; // @[SpriteBlender.scala 81:55]
  wire  _T_2840 = _T_2839 | secondSpriteValids_25; // @[SpriteBlender.scala 81:55]
  wire  _T_2841 = _T_2840 | secondSpriteValids_26; // @[SpriteBlender.scala 81:55]
  wire  _T_2842 = _T_2841 | secondSpriteValids_27; // @[SpriteBlender.scala 81:55]
  wire  _T_2843 = _T_2842 | secondSpriteValids_28; // @[SpriteBlender.scala 81:55]
  wire  _T_2844 = _T_2843 | secondSpriteValids_29; // @[SpriteBlender.scala 81:55]
  wire  _T_2845 = _T_2844 | secondSpriteValids_30; // @[SpriteBlender.scala 81:55]
  wire  _T_2846 = _T_2845 | secondSpriteValids_31; // @[SpriteBlender.scala 81:55]
  wire  _T_2847 = _T_2846 | secondSpriteValids_32; // @[SpriteBlender.scala 81:55]
  wire  _T_2848 = _T_2847 | secondSpriteValids_33; // @[SpriteBlender.scala 81:55]
  wire  _T_2849 = _T_2848 | secondSpriteValids_34; // @[SpriteBlender.scala 81:55]
  wire  _T_2850 = _T_2849 | secondSpriteValids_35; // @[SpriteBlender.scala 81:55]
  wire  _T_2851 = _T_2850 | secondSpriteValids_36; // @[SpriteBlender.scala 81:55]
  wire  _T_2852 = _T_2851 | secondSpriteValids_37; // @[SpriteBlender.scala 81:55]
  wire  _T_2853 = _T_2852 | secondSpriteValids_38; // @[SpriteBlender.scala 81:55]
  wire  _T_2854 = _T_2853 | secondSpriteValids_39; // @[SpriteBlender.scala 81:55]
  wire  _T_2855 = _T_2854 | secondSpriteValids_40; // @[SpriteBlender.scala 81:55]
  wire  _T_2856 = _T_2855 | secondSpriteValids_41; // @[SpriteBlender.scala 81:55]
  wire  _T_2857 = _T_2856 | secondSpriteValids_42; // @[SpriteBlender.scala 81:55]
  wire  _T_2858 = _T_2857 | secondSpriteValids_43; // @[SpriteBlender.scala 81:55]
  wire  _T_2859 = _T_2858 | secondSpriteValids_44; // @[SpriteBlender.scala 81:55]
  wire  _T_2860 = _T_2859 | secondSpriteValids_45; // @[SpriteBlender.scala 81:55]
  wire  _T_2861 = _T_2860 | secondSpriteValids_46; // @[SpriteBlender.scala 81:55]
  wire  _T_2862 = _T_2861 | secondSpriteValids_47; // @[SpriteBlender.scala 81:55]
  wire  _T_2863 = _T_2862 | secondSpriteValids_48; // @[SpriteBlender.scala 81:55]
  wire  _T_2864 = _T_2863 | secondSpriteValids_49; // @[SpriteBlender.scala 81:55]
  wire  _T_2865 = _T_2864 | secondSpriteValids_50; // @[SpriteBlender.scala 81:55]
  wire  _T_2866 = _T_2865 | secondSpriteValids_51; // @[SpriteBlender.scala 81:55]
  wire  _T_2867 = _T_2866 | secondSpriteValids_52; // @[SpriteBlender.scala 81:55]
  wire  _T_2868 = _T_2867 | secondSpriteValids_53; // @[SpriteBlender.scala 81:55]
  wire  _T_2869 = _T_2868 | secondSpriteValids_54; // @[SpriteBlender.scala 81:55]
  wire  _T_2870 = _T_2869 | secondSpriteValids_55; // @[SpriteBlender.scala 81:55]
  wire  _T_2871 = _T_2870 | secondSpriteValids_56; // @[SpriteBlender.scala 81:55]
  wire  _T_2872 = _T_2871 | secondSpriteValids_57; // @[SpriteBlender.scala 81:55]
  wire  _T_2873 = _T_2872 | secondSpriteValids_58; // @[SpriteBlender.scala 81:55]
  wire  _T_2874 = _T_2873 | secondSpriteValids_59; // @[SpriteBlender.scala 81:55]
  wire  _T_2875 = _T_2874 | secondSpriteValids_60; // @[SpriteBlender.scala 81:55]
  wire  _T_2876 = _T_2875 | secondSpriteValids_61; // @[SpriteBlender.scala 81:55]
  wire  _T_2877 = _T_2876 | secondSpriteValids_62; // @[SpriteBlender.scala 81:55]
  wire  _T_2878 = _T_2877 | secondSpriteValids_63; // @[SpriteBlender.scala 81:55]
  wire  _T_2879 = _T_2878 | secondSpriteValids_64; // @[SpriteBlender.scala 81:55]
  wire  _T_2880 = _T_2879 | secondSpriteValids_65; // @[SpriteBlender.scala 81:55]
  wire  _T_2881 = _T_2880 | secondSpriteValids_66; // @[SpriteBlender.scala 81:55]
  wire  _T_2882 = _T_2881 | secondSpriteValids_67; // @[SpriteBlender.scala 81:55]
  wire  _T_2883 = _T_2882 | secondSpriteValids_68; // @[SpriteBlender.scala 81:55]
  wire  _T_2884 = _T_2883 | secondSpriteValids_69; // @[SpriteBlender.scala 81:55]
  wire  _T_2885 = _T_2884 | secondSpriteValids_70; // @[SpriteBlender.scala 81:55]
  wire  _T_2886 = _T_2885 | secondSpriteValids_71; // @[SpriteBlender.scala 81:55]
  wire  _T_2887 = _T_2886 | secondSpriteValids_72; // @[SpriteBlender.scala 81:55]
  wire  _T_2888 = _T_2887 | secondSpriteValids_73; // @[SpriteBlender.scala 81:55]
  wire  _T_2889 = _T_2888 | secondSpriteValids_74; // @[SpriteBlender.scala 81:55]
  wire  _T_2890 = _T_2889 | secondSpriteValids_75; // @[SpriteBlender.scala 81:55]
  wire  _T_2891 = _T_2890 | secondSpriteValids_76; // @[SpriteBlender.scala 81:55]
  wire  _T_2892 = _T_2891 | secondSpriteValids_77; // @[SpriteBlender.scala 81:55]
  wire  _T_2893 = _T_2892 | secondSpriteValids_78; // @[SpriteBlender.scala 81:55]
  wire  _T_2894 = _T_2893 | secondSpriteValids_79; // @[SpriteBlender.scala 81:55]
  wire  _T_2895 = _T_2894 | secondSpriteValids_80; // @[SpriteBlender.scala 81:55]
  wire  _T_2896 = _T_2895 | secondSpriteValids_81; // @[SpriteBlender.scala 81:55]
  wire  _T_2897 = _T_2896 | secondSpriteValids_82; // @[SpriteBlender.scala 81:55]
  wire  _T_2898 = _T_2897 | secondSpriteValids_83; // @[SpriteBlender.scala 81:55]
  wire  _T_2899 = _T_2898 | secondSpriteValids_84; // @[SpriteBlender.scala 81:55]
  wire  _T_2900 = _T_2899 | secondSpriteValids_85; // @[SpriteBlender.scala 81:55]
  wire  _T_2901 = _T_2900 | secondSpriteValids_86; // @[SpriteBlender.scala 81:55]
  wire  _T_2902 = _T_2901 | secondSpriteValids_87; // @[SpriteBlender.scala 81:55]
  wire  _T_2903 = _T_2902 | secondSpriteValids_88; // @[SpriteBlender.scala 81:55]
  wire  _T_2904 = _T_2903 | secondSpriteValids_89; // @[SpriteBlender.scala 81:55]
  wire  _T_2905 = _T_2904 | secondSpriteValids_90; // @[SpriteBlender.scala 81:55]
  wire  _T_2906 = _T_2905 | secondSpriteValids_91; // @[SpriteBlender.scala 81:55]
  wire  _T_2907 = _T_2906 | secondSpriteValids_92; // @[SpriteBlender.scala 81:55]
  wire  _T_2908 = _T_2907 | secondSpriteValids_93; // @[SpriteBlender.scala 81:55]
  wire  _T_2909 = _T_2908 | secondSpriteValids_94; // @[SpriteBlender.scala 81:55]
  wire  _T_2910 = _T_2909 | secondSpriteValids_95; // @[SpriteBlender.scala 81:55]
  wire  _T_2911 = _T_2910 | secondSpriteValids_96; // @[SpriteBlender.scala 81:55]
  wire  _T_2912 = _T_2911 | secondSpriteValids_97; // @[SpriteBlender.scala 81:55]
  wire  _T_2913 = _T_2912 | secondSpriteValids_98; // @[SpriteBlender.scala 81:55]
  wire  _T_2914 = _T_2913 | secondSpriteValids_99; // @[SpriteBlender.scala 81:55]
  wire  _T_2915 = _T_2914 | secondSpriteValids_100; // @[SpriteBlender.scala 81:55]
  wire  _T_2916 = _T_2915 | secondSpriteValids_101; // @[SpriteBlender.scala 81:55]
  wire  _T_2917 = _T_2916 | secondSpriteValids_102; // @[SpriteBlender.scala 81:55]
  wire  _T_2918 = _T_2917 | secondSpriteValids_103; // @[SpriteBlender.scala 81:55]
  wire  _T_2919 = _T_2918 | secondSpriteValids_104; // @[SpriteBlender.scala 81:55]
  wire  _T_2920 = _T_2919 | secondSpriteValids_105; // @[SpriteBlender.scala 81:55]
  wire  _T_2921 = _T_2920 | secondSpriteValids_106; // @[SpriteBlender.scala 81:55]
  wire  _T_2922 = _T_2921 | secondSpriteValids_107; // @[SpriteBlender.scala 81:55]
  wire  _T_2923 = _T_2922 | secondSpriteValids_108; // @[SpriteBlender.scala 81:55]
  wire  _T_2924 = _T_2923 | secondSpriteValids_109; // @[SpriteBlender.scala 81:55]
  wire  _T_2925 = _T_2924 | secondSpriteValids_110; // @[SpriteBlender.scala 81:55]
  wire  _T_2926 = _T_2925 | secondSpriteValids_111; // @[SpriteBlender.scala 81:55]
  wire  _T_2927 = _T_2926 | secondSpriteValids_112; // @[SpriteBlender.scala 81:55]
  wire  _T_2928 = _T_2927 | secondSpriteValids_113; // @[SpriteBlender.scala 81:55]
  wire  _T_2929 = _T_2928 | secondSpriteValids_114; // @[SpriteBlender.scala 81:55]
  wire  _T_2930 = _T_2929 | secondSpriteValids_115; // @[SpriteBlender.scala 81:55]
  wire  _T_2931 = _T_2930 | secondSpriteValids_116; // @[SpriteBlender.scala 81:55]
  wire  _T_2932 = _T_2931 | secondSpriteValids_117; // @[SpriteBlender.scala 81:55]
  wire  _T_2933 = _T_2932 | secondSpriteValids_118; // @[SpriteBlender.scala 81:55]
  wire  _T_2934 = _T_2933 | secondSpriteValids_119; // @[SpriteBlender.scala 81:55]
  wire  _T_2935 = _T_2934 | secondSpriteValids_120; // @[SpriteBlender.scala 81:55]
  wire  _T_2936 = _T_2935 | secondSpriteValids_121; // @[SpriteBlender.scala 81:55]
  wire  _T_2937 = _T_2936 | secondSpriteValids_122; // @[SpriteBlender.scala 81:55]
  wire  _T_2938 = _T_2937 | secondSpriteValids_123; // @[SpriteBlender.scala 81:55]
  wire  _T_2939 = _T_2938 | secondSpriteValids_124; // @[SpriteBlender.scala 81:55]
  wire  _T_2940 = _T_2939 | secondSpriteValids_125; // @[SpriteBlender.scala 81:55]
  wire  _T_2941 = _T_2940 | secondSpriteValids_126; // @[SpriteBlender.scala 81:55]
  wire  secondTopSpriteFound = _T_2941 | secondSpriteValids_127; // @[SpriteBlender.scala 81:55]
  wire  _T_2944 = ~secondTopSpriteFound; // @[SpriteBlender.scala 89:40]
  wire  _T_2950 = secondTopSpriteColor[5:4] > pixelColorBackReg[5:4]; // @[SpriteBlender.scala 95:50]
  wire  _T_2953 = secondTopSpriteColor[3:2] > pixelColorBackReg[3:2]; // @[SpriteBlender.scala 96:50]
  wire  _T_2956 = secondTopSpriteColor[1:0] > pixelColorBackReg[1:0]; // @[SpriteBlender.scala 97:50]
  wire  _T_2959 = ~_T_2950; // @[SpriteBlender.scala 104:40]
  wire  _T_2964 = ~_T_2953; // @[SpriteBlender.scala 106:40]
  wire  _T_2969 = ~_T_2956; // @[SpriteBlender.scala 108:40]
  wire [2:0] _T_2973 = {1'h0,secondTopSpriteColor[5:4]}; // @[SpriteBlender.scala 111:39]
  wire [1:0] _T_2974 = {1'h0,_T_2959}; // @[SpriteBlender.scala 111:65]
  wire [2:0] _GEN_257 = {{1'd0}, _T_2974}; // @[SpriteBlender.scala 111:53]
  wire [2:0] _T_2976 = _T_2973 + _GEN_257; // @[SpriteBlender.scala 111:53]
  wire [2:0] _T_2978 = {1'h0,pixelColorBackReg[5:4]}; // @[SpriteBlender.scala 111:87]
  wire [2:0] _T_2980 = _T_2976 + _T_2978; // @[SpriteBlender.scala 111:75]
  wire [2:0] _T_2983 = {1'h0,secondTopSpriteColor[3:2]}; // @[SpriteBlender.scala 112:39]
  wire [1:0] _T_2984 = {1'h0,_T_2964}; // @[SpriteBlender.scala 112:65]
  wire [2:0] _GEN_258 = {{1'd0}, _T_2984}; // @[SpriteBlender.scala 112:53]
  wire [2:0] _T_2986 = _T_2983 + _GEN_258; // @[SpriteBlender.scala 112:53]
  wire [2:0] _T_2988 = {1'h0,pixelColorBackReg[3:2]}; // @[SpriteBlender.scala 112:87]
  wire [2:0] _T_2990 = _T_2986 + _T_2988; // @[SpriteBlender.scala 112:75]
  wire [2:0] _T_2993 = {1'h0,secondTopSpriteColor[1:0]}; // @[SpriteBlender.scala 113:39]
  wire [1:0] _T_2994 = {1'h0,_T_2969}; // @[SpriteBlender.scala 113:65]
  wire [2:0] _GEN_259 = {{1'd0}, _T_2994}; // @[SpriteBlender.scala 113:53]
  wire [2:0] _T_2996 = _T_2993 + _GEN_259; // @[SpriteBlender.scala 113:53]
  wire [2:0] _T_2998 = {1'h0,pixelColorBackReg[1:0]}; // @[SpriteBlender.scala 113:87]
  wire [2:0] _T_3000 = _T_2996 + _T_2998; // @[SpriteBlender.scala 113:75]
  wire [5:0] _T_3003 = {_T_2980[2:1],_T_2990[2:1],_T_3000[2:1]}; // @[Cat.scala 29:58]
  wire [5:0] blendedColorBot = _T_2944 ? pixelColorBackReg : _T_3003; // @[SpriteBlender.scala 89:63]
  wire  comparerR = topSpriteRGB[5:4] > blendedColorBot[5:4]; // @[SpriteBlender.scala 121:37]
  wire  comparerG = topSpriteRGB[3:2] > blendedColorBot[3:2]; // @[SpriteBlender.scala 122:37]
  wire  comparerB = topSpriteRGB[1:0] > blendedColorBot[1:0]; // @[SpriteBlender.scala 123:37]
  wire  zR = ~comparerR; // @[SpriteBlender.scala 130:35]
  wire  zG = ~comparerG; // @[SpriteBlender.scala 132:35]
  wire  zB = ~comparerB; // @[SpriteBlender.scala 134:35]
  wire [2:0] _T_3025 = {1'h0,topSpriteRGB[5:4]}; // @[SpriteBlender.scala 137:34]
  wire [1:0] _T_3026 = {1'h0,zR}; // @[SpriteBlender.scala 137:56]
  wire [2:0] _GEN_260 = {{1'd0}, _T_3026}; // @[SpriteBlender.scala 137:45]
  wire [2:0] _T_3028 = _T_3025 + _GEN_260; // @[SpriteBlender.scala 137:45]
  wire [2:0] _T_3030 = {1'h0,blendedColorBot[5:4]}; // @[SpriteBlender.scala 137:74]
  wire [2:0] _T_3032 = _T_3028 + _T_3030; // @[SpriteBlender.scala 137:62]
  wire [1:0] blendedColorR = _T_3032[2:1]; // @[SpriteBlender.scala 137:86]
  wire [2:0] _T_3034 = {1'h0,topSpriteRGB[3:2]}; // @[SpriteBlender.scala 138:34]
  wire [1:0] _T_3035 = {1'h0,zG}; // @[SpriteBlender.scala 138:56]
  wire [2:0] _GEN_261 = {{1'd0}, _T_3035}; // @[SpriteBlender.scala 138:45]
  wire [2:0] _T_3037 = _T_3034 + _GEN_261; // @[SpriteBlender.scala 138:45]
  wire [2:0] _T_3039 = {1'h0,blendedColorBot[3:2]}; // @[SpriteBlender.scala 138:74]
  wire [2:0] _T_3041 = _T_3037 + _T_3039; // @[SpriteBlender.scala 138:62]
  wire [1:0] blendedColorG = _T_3041[2:1]; // @[SpriteBlender.scala 138:86]
  wire [2:0] _T_3043 = {1'h0,topSpriteRGB[1:0]}; // @[SpriteBlender.scala 139:34]
  wire [1:0] _T_3044 = {1'h0,zB}; // @[SpriteBlender.scala 139:56]
  wire [2:0] _GEN_262 = {{1'd0}, _T_3044}; // @[SpriteBlender.scala 139:45]
  wire [2:0] _T_3046 = _T_3043 + _GEN_262; // @[SpriteBlender.scala 139:45]
  wire [2:0] _T_3048 = {1'h0,blendedColorBot[1:0]}; // @[SpriteBlender.scala 139:74]
  wire [2:0] _T_3050 = _T_3046 + _T_3048; // @[SpriteBlender.scala 139:62]
  wire [1:0] blendedColorB = _T_3050[2:1]; // @[SpriteBlender.scala 139:86]
  wire  _T_3051 = ~topSpriteAlpha; // @[SpriteBlender.scala 141:44]
  wire  _T_3052 = multiHotPriortyReductionTree_io_selectOutput & _T_3051; // @[SpriteBlender.scala 141:41]
  wire [5:0] _T_3054 = {blendedColorR,blendedColorG,blendedColorB}; // @[Cat.scala 29:58]
  wire [5:0] blendedColor = _T_3052 ? _T_3054 : pixelColorBackReg; // @[SpriteBlender.scala 141:22]
  MultiHotPriortyReductionTree multiHotPriortyReductionTree ( // @[SpriteBlender.scala 33:44]
    .io_dataInput_0(multiHotPriortyReductionTree_io_dataInput_0),
    .io_dataInput_1(multiHotPriortyReductionTree_io_dataInput_1),
    .io_dataInput_2(multiHotPriortyReductionTree_io_dataInput_2),
    .io_dataInput_3(multiHotPriortyReductionTree_io_dataInput_3),
    .io_dataInput_4(multiHotPriortyReductionTree_io_dataInput_4),
    .io_dataInput_5(multiHotPriortyReductionTree_io_dataInput_5),
    .io_dataInput_6(multiHotPriortyReductionTree_io_dataInput_6),
    .io_dataInput_7(multiHotPriortyReductionTree_io_dataInput_7),
    .io_dataInput_8(multiHotPriortyReductionTree_io_dataInput_8),
    .io_dataInput_9(multiHotPriortyReductionTree_io_dataInput_9),
    .io_dataInput_10(multiHotPriortyReductionTree_io_dataInput_10),
    .io_dataInput_11(multiHotPriortyReductionTree_io_dataInput_11),
    .io_dataInput_12(multiHotPriortyReductionTree_io_dataInput_12),
    .io_dataInput_13(multiHotPriortyReductionTree_io_dataInput_13),
    .io_dataInput_14(multiHotPriortyReductionTree_io_dataInput_14),
    .io_dataInput_15(multiHotPriortyReductionTree_io_dataInput_15),
    .io_dataInput_16(multiHotPriortyReductionTree_io_dataInput_16),
    .io_dataInput_17(multiHotPriortyReductionTree_io_dataInput_17),
    .io_dataInput_18(multiHotPriortyReductionTree_io_dataInput_18),
    .io_dataInput_19(multiHotPriortyReductionTree_io_dataInput_19),
    .io_dataInput_20(multiHotPriortyReductionTree_io_dataInput_20),
    .io_dataInput_21(multiHotPriortyReductionTree_io_dataInput_21),
    .io_dataInput_22(multiHotPriortyReductionTree_io_dataInput_22),
    .io_dataInput_23(multiHotPriortyReductionTree_io_dataInput_23),
    .io_dataInput_24(multiHotPriortyReductionTree_io_dataInput_24),
    .io_dataInput_25(multiHotPriortyReductionTree_io_dataInput_25),
    .io_dataInput_26(multiHotPriortyReductionTree_io_dataInput_26),
    .io_dataInput_27(multiHotPriortyReductionTree_io_dataInput_27),
    .io_dataInput_28(multiHotPriortyReductionTree_io_dataInput_28),
    .io_dataInput_29(multiHotPriortyReductionTree_io_dataInput_29),
    .io_dataInput_30(multiHotPriortyReductionTree_io_dataInput_30),
    .io_dataInput_31(multiHotPriortyReductionTree_io_dataInput_31),
    .io_dataInput_32(multiHotPriortyReductionTree_io_dataInput_32),
    .io_dataInput_33(multiHotPriortyReductionTree_io_dataInput_33),
    .io_dataInput_34(multiHotPriortyReductionTree_io_dataInput_34),
    .io_dataInput_35(multiHotPriortyReductionTree_io_dataInput_35),
    .io_dataInput_36(multiHotPriortyReductionTree_io_dataInput_36),
    .io_dataInput_37(multiHotPriortyReductionTree_io_dataInput_37),
    .io_dataInput_38(multiHotPriortyReductionTree_io_dataInput_38),
    .io_dataInput_39(multiHotPriortyReductionTree_io_dataInput_39),
    .io_dataInput_40(multiHotPriortyReductionTree_io_dataInput_40),
    .io_dataInput_41(multiHotPriortyReductionTree_io_dataInput_41),
    .io_dataInput_42(multiHotPriortyReductionTree_io_dataInput_42),
    .io_dataInput_43(multiHotPriortyReductionTree_io_dataInput_43),
    .io_dataInput_44(multiHotPriortyReductionTree_io_dataInput_44),
    .io_dataInput_45(multiHotPriortyReductionTree_io_dataInput_45),
    .io_dataInput_46(multiHotPriortyReductionTree_io_dataInput_46),
    .io_dataInput_47(multiHotPriortyReductionTree_io_dataInput_47),
    .io_dataInput_48(multiHotPriortyReductionTree_io_dataInput_48),
    .io_dataInput_49(multiHotPriortyReductionTree_io_dataInput_49),
    .io_dataInput_50(multiHotPriortyReductionTree_io_dataInput_50),
    .io_dataInput_51(multiHotPriortyReductionTree_io_dataInput_51),
    .io_dataInput_52(multiHotPriortyReductionTree_io_dataInput_52),
    .io_dataInput_53(multiHotPriortyReductionTree_io_dataInput_53),
    .io_dataInput_54(multiHotPriortyReductionTree_io_dataInput_54),
    .io_dataInput_55(multiHotPriortyReductionTree_io_dataInput_55),
    .io_dataInput_56(multiHotPriortyReductionTree_io_dataInput_56),
    .io_dataInput_57(multiHotPriortyReductionTree_io_dataInput_57),
    .io_dataInput_58(multiHotPriortyReductionTree_io_dataInput_58),
    .io_dataInput_59(multiHotPriortyReductionTree_io_dataInput_59),
    .io_dataInput_60(multiHotPriortyReductionTree_io_dataInput_60),
    .io_dataInput_61(multiHotPriortyReductionTree_io_dataInput_61),
    .io_dataInput_62(multiHotPriortyReductionTree_io_dataInput_62),
    .io_dataInput_63(multiHotPriortyReductionTree_io_dataInput_63),
    .io_dataInput_64(multiHotPriortyReductionTree_io_dataInput_64),
    .io_dataInput_65(multiHotPriortyReductionTree_io_dataInput_65),
    .io_dataInput_66(multiHotPriortyReductionTree_io_dataInput_66),
    .io_dataInput_67(multiHotPriortyReductionTree_io_dataInput_67),
    .io_dataInput_68(multiHotPriortyReductionTree_io_dataInput_68),
    .io_dataInput_69(multiHotPriortyReductionTree_io_dataInput_69),
    .io_dataInput_70(multiHotPriortyReductionTree_io_dataInput_70),
    .io_dataInput_71(multiHotPriortyReductionTree_io_dataInput_71),
    .io_dataInput_72(multiHotPriortyReductionTree_io_dataInput_72),
    .io_dataInput_73(multiHotPriortyReductionTree_io_dataInput_73),
    .io_dataInput_74(multiHotPriortyReductionTree_io_dataInput_74),
    .io_dataInput_75(multiHotPriortyReductionTree_io_dataInput_75),
    .io_dataInput_76(multiHotPriortyReductionTree_io_dataInput_76),
    .io_dataInput_77(multiHotPriortyReductionTree_io_dataInput_77),
    .io_dataInput_78(multiHotPriortyReductionTree_io_dataInput_78),
    .io_dataInput_79(multiHotPriortyReductionTree_io_dataInput_79),
    .io_dataInput_80(multiHotPriortyReductionTree_io_dataInput_80),
    .io_dataInput_81(multiHotPriortyReductionTree_io_dataInput_81),
    .io_dataInput_82(multiHotPriortyReductionTree_io_dataInput_82),
    .io_dataInput_83(multiHotPriortyReductionTree_io_dataInput_83),
    .io_dataInput_84(multiHotPriortyReductionTree_io_dataInput_84),
    .io_dataInput_85(multiHotPriortyReductionTree_io_dataInput_85),
    .io_dataInput_86(multiHotPriortyReductionTree_io_dataInput_86),
    .io_dataInput_87(multiHotPriortyReductionTree_io_dataInput_87),
    .io_dataInput_88(multiHotPriortyReductionTree_io_dataInput_88),
    .io_dataInput_89(multiHotPriortyReductionTree_io_dataInput_89),
    .io_dataInput_90(multiHotPriortyReductionTree_io_dataInput_90),
    .io_dataInput_91(multiHotPriortyReductionTree_io_dataInput_91),
    .io_dataInput_92(multiHotPriortyReductionTree_io_dataInput_92),
    .io_dataInput_93(multiHotPriortyReductionTree_io_dataInput_93),
    .io_dataInput_94(multiHotPriortyReductionTree_io_dataInput_94),
    .io_dataInput_95(multiHotPriortyReductionTree_io_dataInput_95),
    .io_dataInput_96(multiHotPriortyReductionTree_io_dataInput_96),
    .io_dataInput_97(multiHotPriortyReductionTree_io_dataInput_97),
    .io_dataInput_98(multiHotPriortyReductionTree_io_dataInput_98),
    .io_dataInput_99(multiHotPriortyReductionTree_io_dataInput_99),
    .io_dataInput_100(multiHotPriortyReductionTree_io_dataInput_100),
    .io_dataInput_101(multiHotPriortyReductionTree_io_dataInput_101),
    .io_dataInput_102(multiHotPriortyReductionTree_io_dataInput_102),
    .io_dataInput_103(multiHotPriortyReductionTree_io_dataInput_103),
    .io_dataInput_104(multiHotPriortyReductionTree_io_dataInput_104),
    .io_dataInput_105(multiHotPriortyReductionTree_io_dataInput_105),
    .io_dataInput_106(multiHotPriortyReductionTree_io_dataInput_106),
    .io_dataInput_107(multiHotPriortyReductionTree_io_dataInput_107),
    .io_dataInput_108(multiHotPriortyReductionTree_io_dataInput_108),
    .io_dataInput_109(multiHotPriortyReductionTree_io_dataInput_109),
    .io_dataInput_110(multiHotPriortyReductionTree_io_dataInput_110),
    .io_dataInput_111(multiHotPriortyReductionTree_io_dataInput_111),
    .io_dataInput_112(multiHotPriortyReductionTree_io_dataInput_112),
    .io_dataInput_113(multiHotPriortyReductionTree_io_dataInput_113),
    .io_dataInput_114(multiHotPriortyReductionTree_io_dataInput_114),
    .io_dataInput_115(multiHotPriortyReductionTree_io_dataInput_115),
    .io_dataInput_116(multiHotPriortyReductionTree_io_dataInput_116),
    .io_dataInput_117(multiHotPriortyReductionTree_io_dataInput_117),
    .io_dataInput_118(multiHotPriortyReductionTree_io_dataInput_118),
    .io_dataInput_119(multiHotPriortyReductionTree_io_dataInput_119),
    .io_dataInput_120(multiHotPriortyReductionTree_io_dataInput_120),
    .io_dataInput_121(multiHotPriortyReductionTree_io_dataInput_121),
    .io_dataInput_122(multiHotPriortyReductionTree_io_dataInput_122),
    .io_dataInput_123(multiHotPriortyReductionTree_io_dataInput_123),
    .io_dataInput_124(multiHotPriortyReductionTree_io_dataInput_124),
    .io_dataInput_125(multiHotPriortyReductionTree_io_dataInput_125),
    .io_dataInput_126(multiHotPriortyReductionTree_io_dataInput_126),
    .io_dataInput_127(multiHotPriortyReductionTree_io_dataInput_127),
    .io_selectInput_0(multiHotPriortyReductionTree_io_selectInput_0),
    .io_selectInput_1(multiHotPriortyReductionTree_io_selectInput_1),
    .io_selectInput_2(multiHotPriortyReductionTree_io_selectInput_2),
    .io_selectInput_3(multiHotPriortyReductionTree_io_selectInput_3),
    .io_selectInput_4(multiHotPriortyReductionTree_io_selectInput_4),
    .io_selectInput_5(multiHotPriortyReductionTree_io_selectInput_5),
    .io_selectInput_6(multiHotPriortyReductionTree_io_selectInput_6),
    .io_selectInput_7(multiHotPriortyReductionTree_io_selectInput_7),
    .io_selectInput_8(multiHotPriortyReductionTree_io_selectInput_8),
    .io_selectInput_9(multiHotPriortyReductionTree_io_selectInput_9),
    .io_selectInput_10(multiHotPriortyReductionTree_io_selectInput_10),
    .io_selectInput_11(multiHotPriortyReductionTree_io_selectInput_11),
    .io_selectInput_12(multiHotPriortyReductionTree_io_selectInput_12),
    .io_selectInput_13(multiHotPriortyReductionTree_io_selectInput_13),
    .io_selectInput_14(multiHotPriortyReductionTree_io_selectInput_14),
    .io_selectInput_15(multiHotPriortyReductionTree_io_selectInput_15),
    .io_selectInput_16(multiHotPriortyReductionTree_io_selectInput_16),
    .io_selectInput_17(multiHotPriortyReductionTree_io_selectInput_17),
    .io_selectInput_18(multiHotPriortyReductionTree_io_selectInput_18),
    .io_selectInput_19(multiHotPriortyReductionTree_io_selectInput_19),
    .io_selectInput_20(multiHotPriortyReductionTree_io_selectInput_20),
    .io_selectInput_21(multiHotPriortyReductionTree_io_selectInput_21),
    .io_selectInput_22(multiHotPriortyReductionTree_io_selectInput_22),
    .io_selectInput_23(multiHotPriortyReductionTree_io_selectInput_23),
    .io_selectInput_24(multiHotPriortyReductionTree_io_selectInput_24),
    .io_selectInput_25(multiHotPriortyReductionTree_io_selectInput_25),
    .io_selectInput_26(multiHotPriortyReductionTree_io_selectInput_26),
    .io_selectInput_27(multiHotPriortyReductionTree_io_selectInput_27),
    .io_selectInput_28(multiHotPriortyReductionTree_io_selectInput_28),
    .io_selectInput_29(multiHotPriortyReductionTree_io_selectInput_29),
    .io_selectInput_30(multiHotPriortyReductionTree_io_selectInput_30),
    .io_selectInput_31(multiHotPriortyReductionTree_io_selectInput_31),
    .io_selectInput_32(multiHotPriortyReductionTree_io_selectInput_32),
    .io_selectInput_33(multiHotPriortyReductionTree_io_selectInput_33),
    .io_selectInput_34(multiHotPriortyReductionTree_io_selectInput_34),
    .io_selectInput_35(multiHotPriortyReductionTree_io_selectInput_35),
    .io_selectInput_36(multiHotPriortyReductionTree_io_selectInput_36),
    .io_selectInput_37(multiHotPriortyReductionTree_io_selectInput_37),
    .io_selectInput_38(multiHotPriortyReductionTree_io_selectInput_38),
    .io_selectInput_39(multiHotPriortyReductionTree_io_selectInput_39),
    .io_selectInput_40(multiHotPriortyReductionTree_io_selectInput_40),
    .io_selectInput_41(multiHotPriortyReductionTree_io_selectInput_41),
    .io_selectInput_42(multiHotPriortyReductionTree_io_selectInput_42),
    .io_selectInput_43(multiHotPriortyReductionTree_io_selectInput_43),
    .io_selectInput_44(multiHotPriortyReductionTree_io_selectInput_44),
    .io_selectInput_45(multiHotPriortyReductionTree_io_selectInput_45),
    .io_selectInput_46(multiHotPriortyReductionTree_io_selectInput_46),
    .io_selectInput_47(multiHotPriortyReductionTree_io_selectInput_47),
    .io_selectInput_48(multiHotPriortyReductionTree_io_selectInput_48),
    .io_selectInput_49(multiHotPriortyReductionTree_io_selectInput_49),
    .io_selectInput_50(multiHotPriortyReductionTree_io_selectInput_50),
    .io_selectInput_51(multiHotPriortyReductionTree_io_selectInput_51),
    .io_selectInput_52(multiHotPriortyReductionTree_io_selectInput_52),
    .io_selectInput_53(multiHotPriortyReductionTree_io_selectInput_53),
    .io_selectInput_54(multiHotPriortyReductionTree_io_selectInput_54),
    .io_selectInput_55(multiHotPriortyReductionTree_io_selectInput_55),
    .io_selectInput_56(multiHotPriortyReductionTree_io_selectInput_56),
    .io_selectInput_57(multiHotPriortyReductionTree_io_selectInput_57),
    .io_selectInput_58(multiHotPriortyReductionTree_io_selectInput_58),
    .io_selectInput_59(multiHotPriortyReductionTree_io_selectInput_59),
    .io_selectInput_60(multiHotPriortyReductionTree_io_selectInput_60),
    .io_selectInput_61(multiHotPriortyReductionTree_io_selectInput_61),
    .io_selectInput_62(multiHotPriortyReductionTree_io_selectInput_62),
    .io_selectInput_63(multiHotPriortyReductionTree_io_selectInput_63),
    .io_selectInput_64(multiHotPriortyReductionTree_io_selectInput_64),
    .io_selectInput_65(multiHotPriortyReductionTree_io_selectInput_65),
    .io_selectInput_66(multiHotPriortyReductionTree_io_selectInput_66),
    .io_selectInput_67(multiHotPriortyReductionTree_io_selectInput_67),
    .io_selectInput_68(multiHotPriortyReductionTree_io_selectInput_68),
    .io_selectInput_69(multiHotPriortyReductionTree_io_selectInput_69),
    .io_selectInput_70(multiHotPriortyReductionTree_io_selectInput_70),
    .io_selectInput_71(multiHotPriortyReductionTree_io_selectInput_71),
    .io_selectInput_72(multiHotPriortyReductionTree_io_selectInput_72),
    .io_selectInput_73(multiHotPriortyReductionTree_io_selectInput_73),
    .io_selectInput_74(multiHotPriortyReductionTree_io_selectInput_74),
    .io_selectInput_75(multiHotPriortyReductionTree_io_selectInput_75),
    .io_selectInput_76(multiHotPriortyReductionTree_io_selectInput_76),
    .io_selectInput_77(multiHotPriortyReductionTree_io_selectInput_77),
    .io_selectInput_78(multiHotPriortyReductionTree_io_selectInput_78),
    .io_selectInput_79(multiHotPriortyReductionTree_io_selectInput_79),
    .io_selectInput_80(multiHotPriortyReductionTree_io_selectInput_80),
    .io_selectInput_81(multiHotPriortyReductionTree_io_selectInput_81),
    .io_selectInput_82(multiHotPriortyReductionTree_io_selectInput_82),
    .io_selectInput_83(multiHotPriortyReductionTree_io_selectInput_83),
    .io_selectInput_84(multiHotPriortyReductionTree_io_selectInput_84),
    .io_selectInput_85(multiHotPriortyReductionTree_io_selectInput_85),
    .io_selectInput_86(multiHotPriortyReductionTree_io_selectInput_86),
    .io_selectInput_87(multiHotPriortyReductionTree_io_selectInput_87),
    .io_selectInput_88(multiHotPriortyReductionTree_io_selectInput_88),
    .io_selectInput_89(multiHotPriortyReductionTree_io_selectInput_89),
    .io_selectInput_90(multiHotPriortyReductionTree_io_selectInput_90),
    .io_selectInput_91(multiHotPriortyReductionTree_io_selectInput_91),
    .io_selectInput_92(multiHotPriortyReductionTree_io_selectInput_92),
    .io_selectInput_93(multiHotPriortyReductionTree_io_selectInput_93),
    .io_selectInput_94(multiHotPriortyReductionTree_io_selectInput_94),
    .io_selectInput_95(multiHotPriortyReductionTree_io_selectInput_95),
    .io_selectInput_96(multiHotPriortyReductionTree_io_selectInput_96),
    .io_selectInput_97(multiHotPriortyReductionTree_io_selectInput_97),
    .io_selectInput_98(multiHotPriortyReductionTree_io_selectInput_98),
    .io_selectInput_99(multiHotPriortyReductionTree_io_selectInput_99),
    .io_selectInput_100(multiHotPriortyReductionTree_io_selectInput_100),
    .io_selectInput_101(multiHotPriortyReductionTree_io_selectInput_101),
    .io_selectInput_102(multiHotPriortyReductionTree_io_selectInput_102),
    .io_selectInput_103(multiHotPriortyReductionTree_io_selectInput_103),
    .io_selectInput_104(multiHotPriortyReductionTree_io_selectInput_104),
    .io_selectInput_105(multiHotPriortyReductionTree_io_selectInput_105),
    .io_selectInput_106(multiHotPriortyReductionTree_io_selectInput_106),
    .io_selectInput_107(multiHotPriortyReductionTree_io_selectInput_107),
    .io_selectInput_108(multiHotPriortyReductionTree_io_selectInput_108),
    .io_selectInput_109(multiHotPriortyReductionTree_io_selectInput_109),
    .io_selectInput_110(multiHotPriortyReductionTree_io_selectInput_110),
    .io_selectInput_111(multiHotPriortyReductionTree_io_selectInput_111),
    .io_selectInput_112(multiHotPriortyReductionTree_io_selectInput_112),
    .io_selectInput_113(multiHotPriortyReductionTree_io_selectInput_113),
    .io_selectInput_114(multiHotPriortyReductionTree_io_selectInput_114),
    .io_selectInput_115(multiHotPriortyReductionTree_io_selectInput_115),
    .io_selectInput_116(multiHotPriortyReductionTree_io_selectInput_116),
    .io_selectInput_117(multiHotPriortyReductionTree_io_selectInput_117),
    .io_selectInput_118(multiHotPriortyReductionTree_io_selectInput_118),
    .io_selectInput_119(multiHotPriortyReductionTree_io_selectInput_119),
    .io_selectInput_120(multiHotPriortyReductionTree_io_selectInput_120),
    .io_selectInput_121(multiHotPriortyReductionTree_io_selectInput_121),
    .io_selectInput_122(multiHotPriortyReductionTree_io_selectInput_122),
    .io_selectInput_123(multiHotPriortyReductionTree_io_selectInput_123),
    .io_selectInput_124(multiHotPriortyReductionTree_io_selectInput_124),
    .io_selectInput_125(multiHotPriortyReductionTree_io_selectInput_125),
    .io_selectInput_126(multiHotPriortyReductionTree_io_selectInput_126),
    .io_selectInput_127(multiHotPriortyReductionTree_io_selectInput_127),
    .io_dataOutput(multiHotPriortyReductionTree_io_dataOutput),
    .io_selectOutput(multiHotPriortyReductionTree_io_selectOutput),
    .io_indexOutput(multiHotPriortyReductionTree_io_indexOutput)
  );
  assign io_vgaRed = {blendedColor[5:4],blendedColor[5:4]}; // @[SpriteBlender.scala 152:13 SpriteBlender.scala 157:13]
  assign io_vgaGreen = {blendedColor[3:2],blendedColor[3:2]}; // @[SpriteBlender.scala 153:15 SpriteBlender.scala 158:15]
  assign io_vgaBlue = {blendedColor[1:0],blendedColor[1:0]}; // @[SpriteBlender.scala 154:14 SpriteBlender.scala 159:14]
  assign multiHotPriortyReductionTree_io_dataInput_0 = io_datareader_0; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_1 = io_datareader_1; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_2 = io_datareader_2; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_3 = io_datareader_3; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_4 = io_datareader_4; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_5 = io_datareader_5; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_6 = io_datareader_6; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_7 = io_datareader_7; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_8 = io_datareader_8; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_9 = io_datareader_9; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_10 = io_datareader_10; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_11 = io_datareader_11; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_12 = io_datareader_12; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_13 = io_datareader_13; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_14 = io_datareader_14; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_15 = io_datareader_15; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_16 = io_datareader_16; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_17 = io_datareader_17; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_18 = io_datareader_18; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_19 = io_datareader_19; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_20 = io_datareader_20; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_21 = io_datareader_21; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_22 = io_datareader_22; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_23 = io_datareader_23; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_24 = io_datareader_24; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_25 = io_datareader_25; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_26 = io_datareader_26; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_27 = io_datareader_27; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_28 = io_datareader_28; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_29 = io_datareader_29; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_30 = io_datareader_30; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_31 = io_datareader_31; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_32 = io_datareader_32; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_33 = io_datareader_33; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_34 = io_datareader_34; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_35 = io_datareader_35; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_36 = io_datareader_36; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_37 = io_datareader_37; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_38 = io_datareader_38; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_39 = io_datareader_39; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_40 = io_datareader_40; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_41 = io_datareader_41; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_42 = io_datareader_42; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_43 = io_datareader_43; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_44 = io_datareader_44; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_45 = io_datareader_45; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_46 = io_datareader_46; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_47 = io_datareader_47; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_48 = io_datareader_48; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_49 = io_datareader_49; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_50 = io_datareader_50; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_51 = io_datareader_51; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_52 = io_datareader_52; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_53 = io_datareader_53; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_54 = io_datareader_54; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_55 = io_datareader_55; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_56 = io_datareader_56; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_57 = io_datareader_57; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_58 = io_datareader_58; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_59 = io_datareader_59; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_60 = io_datareader_60; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_61 = io_datareader_61; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_62 = io_datareader_62; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_63 = io_datareader_63; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_64 = io_datareader_64; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_65 = io_datareader_65; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_66 = io_datareader_66; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_67 = io_datareader_67; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_68 = io_datareader_68; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_69 = io_datareader_69; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_70 = io_datareader_70; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_71 = io_datareader_71; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_72 = io_datareader_72; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_73 = io_datareader_73; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_74 = io_datareader_74; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_75 = io_datareader_75; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_76 = io_datareader_76; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_77 = io_datareader_77; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_78 = io_datareader_78; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_79 = io_datareader_79; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_80 = io_datareader_80; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_81 = io_datareader_81; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_82 = io_datareader_82; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_83 = io_datareader_83; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_84 = io_datareader_84; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_85 = io_datareader_85; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_86 = io_datareader_86; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_87 = io_datareader_87; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_88 = io_datareader_88; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_89 = io_datareader_89; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_90 = io_datareader_90; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_91 = io_datareader_91; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_92 = io_datareader_92; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_93 = io_datareader_93; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_94 = io_datareader_94; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_95 = io_datareader_95; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_96 = io_datareader_96; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_97 = io_datareader_97; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_98 = io_datareader_98; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_99 = io_datareader_99; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_100 = io_datareader_100; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_101 = io_datareader_101; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_102 = io_datareader_102; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_103 = io_datareader_103; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_104 = io_datareader_104; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_105 = io_datareader_105; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_106 = io_datareader_106; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_107 = io_datareader_107; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_108 = io_datareader_108; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_109 = io_datareader_109; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_110 = io_datareader_110; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_111 = io_datareader_111; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_112 = io_datareader_112; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_113 = io_datareader_113; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_114 = io_datareader_114; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_115 = io_datareader_115; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_116 = io_datareader_116; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_117 = io_datareader_117; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_118 = io_datareader_118; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_119 = io_datareader_119; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_120 = io_datareader_120; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_121 = io_datareader_121; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_122 = io_datareader_122; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_123 = io_datareader_123; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_124 = io_datareader_124; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_125 = io_datareader_125; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_126 = io_datareader_126; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_dataInput_127 = io_datareader_127; // @[SpriteBlender.scala 36:50]
  assign multiHotPriortyReductionTree_io_selectInput_0 = _T_5 & _T_7; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_1 = _T_13 & _T_15; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_2 = _T_21 & _T_23; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_3 = _T_29 & _T_31; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_4 = _T_37 & _T_39; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_5 = _T_45 & _T_47; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_6 = _T_53 & _T_55; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_7 = _T_61 & _T_63; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_8 = _T_69 & _T_71; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_9 = _T_77 & _T_79; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_10 = _T_85 & _T_87; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_11 = _T_93 & _T_95; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_12 = _T_101 & _T_103; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_13 = _T_109 & _T_111; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_14 = _T_117 & _T_119; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_15 = _T_125 & _T_127; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_16 = _T_133 & _T_135; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_17 = _T_141 & _T_143; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_18 = _T_149 & _T_151; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_19 = _T_157 & _T_159; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_20 = _T_165 & _T_167; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_21 = _T_173 & _T_175; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_22 = _T_181 & _T_183; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_23 = _T_189 & _T_191; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_24 = _T_197 & _T_199; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_25 = _T_205 & _T_207; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_26 = _T_213 & _T_215; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_27 = _T_221 & _T_223; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_28 = _T_229 & _T_231; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_29 = _T_237 & _T_239; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_30 = _T_245 & _T_247; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_31 = _T_253 & _T_255; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_32 = _T_261 & _T_263; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_33 = _T_269 & _T_271; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_34 = _T_276_0 & _T_279; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_35 = _T_284_0 & _T_287; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_36 = _T_292_0 & _T_295; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_37 = _T_300_0 & _T_303; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_38 = _T_308_0 & _T_311; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_39 = _T_316_0 & _T_319; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_40 = _T_324_0 & _T_327; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_41 = _T_333 & _T_335; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_42 = _T_341 & _T_343; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_43 = _T_349 & _T_351; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_44 = _T_357 & _T_359; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_45 = _T_365 & _T_367; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_46 = _T_373 & _T_375; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_47 = _T_381 & _T_383; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_48 = _T_389 & _T_391; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_49 = _T_397 & _T_399; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_50 = _T_405 & _T_407; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_51 = _T_413 & _T_415; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_52 = _T_420_0 & _T_423; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_53 = _T_428_0 & _T_431; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_54 = _T_436_0 & _T_439; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_55 = _T_445 & _T_447; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_56 = _T_453 & _T_455; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_57 = _T_461 & _T_463; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_58 = _T_468_0 & _T_471; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_59 = _T_476_0 & _T_479; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_60 = _T_484_0 & _T_487; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_61 = _T_493 & _T_495; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_62 = _T_501 & _T_503; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_63 = _T_509 & _T_511; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_64 = _T_517 & _T_519; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_65 = _T_525 & _T_527; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_66 = _T_533 & _T_535; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_67 = _T_540_0 & _T_543; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_68 = _T_548_0 & _T_551; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_69 = _T_556_0 & _T_559; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_70 = _T_565 & _T_567; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_71 = _T_573 & _T_575; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_72 = _T_581 & _T_583; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_73 = _T_588_0 & _T_591; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_74 = _T_596_0 & _T_599; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_75 = _T_604_0 & _T_607; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_76 = _T_612_0 & _T_615; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_77 = _T_620_0 & _T_623; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_78 = _T_628_0 & _T_631; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_79 = _T_636_0 & _T_639; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_80 = _T_644_0 & _T_647; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_81 = _T_652_0 & _T_655; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_82 = _T_660_0 & _T_663; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_83 = _T_668_0 & _T_671; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_84 = _T_676_0 & _T_679; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_85 = _T_684_0 & _T_687; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_86 = _T_692_0 & _T_695; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_87 = _T_700_0 & _T_703; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_88 = _T_708_0 & _T_711; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_89 = _T_716_0 & _T_719; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_90 = _T_724_0 & _T_727; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_91 = _T_732_0 & _T_735; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_92 = _T_740_0 & _T_743; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_93 = _T_748_0 & _T_751; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_94 = _T_756_0 & _T_759; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_95 = _T_764_0 & _T_767; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_96 = _T_772_0 & _T_775; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_97 = _T_780_0 & _T_783; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_98 = _T_788_0 & _T_791; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_99 = _T_796_0 & _T_799; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_100 = _T_804_0 & _T_807; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_101 = _T_812_0 & _T_815; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_102 = _T_820_0 & _T_823; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_103 = _T_828_0 & _T_831; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_104 = _T_836_0 & _T_839; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_105 = _T_844_0 & _T_847; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_106 = _T_852_0 & _T_855; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_107 = _T_860_0 & _T_863; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_108 = _T_868_0 & _T_871; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_109 = _T_876_0 & _T_879; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_110 = _T_884_0 & _T_887; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_111 = _T_892_0 & _T_895; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_112 = _T_900_0 & _T_903; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_113 = _T_908_0 & _T_911; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_114 = _T_916_0 & _T_919; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_115 = _T_924_0 & _T_927; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_116 = _T_932_0 & _T_935; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_117 = _T_940_0 & _T_943; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_118 = _T_948_0 & _T_951; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_119 = _T_956_0 & _T_959; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_120 = _T_964_0 & _T_967; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_121 = _T_972_0 & _T_975; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_122 = _T_980_0 & _T_983; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_123 = _T_988_0 & _T_991; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_124 = _T_996_0 & _T_999; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_125 = _T_1004_0 & _T_1007; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_126 = _T_1012_0 & _T_1015; // @[SpriteBlender.scala 39:52]
  assign multiHotPriortyReductionTree_io_selectInput_127 = _T_1020_0 & _T_1023; // @[SpriteBlender.scala 39:52]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  pixelColorBackReg = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_3_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_4_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_4_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_11_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_11_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_12_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_12_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_19_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_19_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_20_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_20_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_27_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_27_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_28_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_28_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_35_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_35_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_36_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_36_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_43_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_43_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_44_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_44_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_51_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_51_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_52_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_52_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_59_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_59_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_60_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_60_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_67_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_67_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_68_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_68_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_75_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_75_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_76_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_76_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_83_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_83_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_84_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_84_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_91_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_91_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_92_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_92_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_99_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_99_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_100_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_100_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _T_107_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _T_107_1 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_108_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_108_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _T_115_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _T_115_1 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  _T_116_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_116_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_123_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_123_1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_124_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_124_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _T_131_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  _T_131_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _T_132_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _T_132_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _T_139_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _T_139_1 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _T_140_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _T_140_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _T_147_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  _T_147_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _T_148_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  _T_148_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  _T_155_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  _T_155_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  _T_156_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  _T_156_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  _T_163_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  _T_163_1 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  _T_164_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  _T_164_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  _T_171_0 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _T_171_1 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _T_172_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  _T_172_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _T_179_0 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  _T_179_1 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  _T_180_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _T_180_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_187_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _T_187_1 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _T_188_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _T_188_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _T_195_0 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _T_195_1 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _T_196_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  _T_196_1 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  _T_203_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  _T_203_1 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  _T_204_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _T_204_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  _T_211_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  _T_211_1 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _T_212_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  _T_212_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  _T_219_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  _T_219_1 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  _T_220_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  _T_220_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  _T_227_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  _T_227_1 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  _T_228_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  _T_228_1 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  _T_235_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  _T_235_1 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  _T_236_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  _T_236_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  _T_243_0 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  _T_243_1 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  _T_244_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  _T_244_1 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  _T_251_0 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  _T_251_1 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  _T_252_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  _T_252_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  _T_259_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  _T_259_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  _T_260_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _T_260_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  _T_267_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  _T_267_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _T_268_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  _T_268_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _T_276_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  _T_276_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  _T_284_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  _T_284_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _T_292_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  _T_292_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _T_300_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  _T_300_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  _T_308_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _T_308_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _T_316_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  _T_316_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _T_324_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  _T_324_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  _T_331_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  _T_331_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _T_332_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  _T_332_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _T_339_0 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _T_339_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _T_340_0 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  _T_340_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _T_347_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  _T_347_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _T_348_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  _T_348_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  _T_355_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _T_355_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _T_356_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_356_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  _T_363_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  _T_363_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  _T_364_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  _T_364_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _T_371_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  _T_371_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_372_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  _T_372_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  _T_379_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_379_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _T_380_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _T_380_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _T_387_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  _T_387_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  _T_388_0 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  _T_388_1 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  _T_395_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  _T_395_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  _T_396_0 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  _T_396_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  _T_403_0 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  _T_403_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  _T_404_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  _T_404_1 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  _T_411_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  _T_411_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  _T_412_0 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  _T_412_1 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  _T_420_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  _T_420_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  _T_428_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  _T_428_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  _T_436_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  _T_436_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  _T_443_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  _T_443_1 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  _T_444_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  _T_444_1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  _T_451_0 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  _T_451_1 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  _T_452_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  _T_452_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  _T_459_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  _T_459_1 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  _T_460_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  _T_460_1 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  _T_468_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  _T_468_1 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  _T_476_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  _T_476_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  _T_484_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  _T_484_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  _T_491_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  _T_491_1 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  _T_492_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  _T_492_1 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  _T_499_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  _T_499_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  _T_500_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  _T_500_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  _T_507_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  _T_507_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  _T_508_0 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  _T_508_1 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  _T_515_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  _T_515_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  _T_516_0 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  _T_516_1 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  _T_523_0 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  _T_523_1 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  _T_524_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  _T_524_1 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  _T_531_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  _T_531_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  _T_532_0 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  _T_532_1 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  _T_540_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  _T_540_1 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  _T_548_0 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  _T_548_1 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  _T_556_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  _T_556_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  _T_563_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  _T_563_1 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  _T_564_0 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  _T_564_1 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  _T_571_0 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  _T_571_1 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  _T_572_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  _T_572_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  _T_579_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  _T_579_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  _T_580_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  _T_580_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  _T_588_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  _T_588_1 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  _T_596_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  _T_596_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  _T_604_0 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  _T_604_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  _T_612_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  _T_612_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  _T_620_0 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  _T_620_1 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  _T_628_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  _T_628_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  _T_636_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  _T_636_1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  _T_644_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  _T_644_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_652_0 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  _T_652_1 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  _T_660_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  _T_660_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  _T_668_0 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  _T_668_1 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_676_0 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  _T_676_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  _T_684_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  _T_684_1 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  _T_692_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  _T_692_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  _T_700_0 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  _T_700_1 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  _T_708_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  _T_708_1 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  _T_716_0 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  _T_716_1 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  _T_724_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  _T_724_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  _T_732_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  _T_732_1 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  _T_740_0 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  _T_740_1 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  _T_748_0 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  _T_748_1 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  _T_756_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  _T_756_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  _T_764_0 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  _T_764_1 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  _T_772_0 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  _T_772_1 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  _T_780_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  _T_780_1 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  _T_788_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  _T_788_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  _T_796_0 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  _T_796_1 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  _T_804_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  _T_804_1 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  _T_812_0 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  _T_812_1 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  _T_820_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  _T_820_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  _T_828_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  _T_828_1 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  _T_836_0 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  _T_836_1 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  _T_844_0 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  _T_844_1 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  _T_852_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  _T_852_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  _T_860_0 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  _T_860_1 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  _T_868_0 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  _T_868_1 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  _T_876_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  _T_876_1 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  _T_884_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  _T_884_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  _T_892_0 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  _T_892_1 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  _T_900_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  _T_900_1 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  _T_908_0 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  _T_908_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  _T_916_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  _T_916_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  _T_924_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  _T_924_1 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  _T_932_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  _T_932_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  _T_940_0 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  _T_940_1 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  _T_948_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  _T_948_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  _T_956_0 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  _T_956_1 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  _T_964_0 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  _T_964_1 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  _T_972_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  _T_972_1 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  _T_980_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  _T_980_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  _T_988_0 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  _T_988_1 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  _T_996_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  _T_996_1 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  _T_1004_0 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  _T_1004_1 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  _T_1012_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  _T_1012_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  _T_1020_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  _T_1020_1 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  _T_1026_0 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  _T_1026_1 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  _T_1027_0 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  _T_1027_1 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  _T_1038_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  _T_1038_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  _T_1039_0 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  _T_1039_1 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  _T_1050_0 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  _T_1050_1 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  _T_1051_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  _T_1051_1 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  _T_1062_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  _T_1062_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  _T_1063_0 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  _T_1063_1 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  _T_1074_0 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  _T_1074_1 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  _T_1075_0 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  _T_1075_1 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  _T_1086_0 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  _T_1086_1 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  _T_1087_0 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  _T_1087_1 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  _T_1098_0 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  _T_1098_1 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  _T_1099_0 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  _T_1099_1 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  _T_1110_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  _T_1110_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  _T_1111_0 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  _T_1111_1 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  _T_1122_0 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  _T_1122_1 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  _T_1123_0 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  _T_1123_1 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  _T_1134_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  _T_1134_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  _T_1135_0 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  _T_1135_1 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  _T_1146_0 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  _T_1146_1 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  _T_1147_0 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  _T_1147_1 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  _T_1158_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  _T_1158_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  _T_1159_0 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  _T_1159_1 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  _T_1170_0 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  _T_1170_1 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  _T_1171_0 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  _T_1171_1 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  _T_1182_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  _T_1182_1 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  _T_1183_0 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  _T_1183_1 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  _T_1194_0 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  _T_1194_1 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  _T_1195_0 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  _T_1195_1 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  _T_1206_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  _T_1206_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  _T_1207_0 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  _T_1207_1 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  _T_1218_0 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  _T_1218_1 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  _T_1219_0 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  _T_1219_1 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  _T_1230_0 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  _T_1230_1 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  _T_1231_0 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  _T_1231_1 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  _T_1242_0 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  _T_1242_1 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  _T_1243_0 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  _T_1243_1 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  _T_1254_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  _T_1254_1 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  _T_1255_0 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  _T_1255_1 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  _T_1266_0 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  _T_1266_1 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  _T_1267_0 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  _T_1267_1 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  _T_1278_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  _T_1278_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  _T_1279_0 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  _T_1279_1 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  _T_1290_0 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  _T_1290_1 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  _T_1291_0 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_1291_1 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_1302_0 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_1302_1 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_1303_0 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_1303_1 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_1314_0 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_1314_1 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_1315_0 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_1315_1 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_1326_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  _T_1326_1 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  _T_1327_0 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  _T_1327_1 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  _T_1338_0 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  _T_1338_1 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  _T_1339_0 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  _T_1339_1 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  _T_1350_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  _T_1350_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  _T_1351_0 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  _T_1351_1 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  _T_1362_0 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  _T_1362_1 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  _T_1363_0 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  _T_1363_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  _T_1374_0 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  _T_1374_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  _T_1375_0 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  _T_1375_1 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  _T_1386_0 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  _T_1386_1 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  _T_1387_0 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  _T_1387_1 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  _T_1398_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  _T_1398_1 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  _T_1399_0 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  _T_1399_1 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  _T_1410_0 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  _T_1410_1 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  _T_1411_0 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  _T_1411_1 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  _T_1422_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  _T_1422_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  _T_1423_0 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  _T_1423_1 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  _T_1435_0 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  _T_1435_1 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  _T_1447_0 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  _T_1447_1 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  _T_1459_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  _T_1459_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  _T_1471_0 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  _T_1471_1 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  _T_1483_0 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  _T_1483_1 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  _T_1495_0 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  _T_1495_1 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  _T_1507_0 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  _T_1507_1 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  _T_1518_0 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  _T_1518_1 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  _T_1519_0 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  _T_1519_1 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  _T_1530_0 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  _T_1530_1 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  _T_1531_0 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  _T_1531_1 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  _T_1542_0 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  _T_1542_1 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  _T_1543_0 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  _T_1543_1 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  _T_1554_0 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  _T_1554_1 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  _T_1555_0 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  _T_1555_1 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  _T_1566_0 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  _T_1566_1 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  _T_1567_0 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  _T_1567_1 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  _T_1578_0 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  _T_1578_1 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  _T_1579_0 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  _T_1579_1 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  _T_1590_0 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  _T_1590_1 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  _T_1591_0 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  _T_1591_1 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  _T_1602_0 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  _T_1602_1 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  _T_1603_0 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  _T_1603_1 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  _T_1614_0 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  _T_1614_1 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  _T_1615_0 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  _T_1615_1 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  _T_1626_0 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  _T_1626_1 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  _T_1627_0 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  _T_1627_1 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  _T_1638_0 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  _T_1638_1 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  _T_1639_0 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  _T_1639_1 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  _T_1651_0 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  _T_1651_1 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  _T_1663_0 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  _T_1663_1 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  _T_1675_0 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  _T_1675_1 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  _T_1686_0 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  _T_1686_1 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  _T_1687_0 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  _T_1687_1 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  _T_1698_0 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  _T_1698_1 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  _T_1699_0 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  _T_1699_1 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  _T_1710_0 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  _T_1710_1 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  _T_1711_0 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  _T_1711_1 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  _T_1723_0 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  _T_1723_1 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  _T_1735_0 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  _T_1735_1 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  _T_1747_0 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  _T_1747_1 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  _T_1758_0 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  _T_1758_1 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  _T_1759_0 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  _T_1759_1 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  _T_1770_0 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  _T_1770_1 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  _T_1771_0 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  _T_1771_1 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  _T_1782_0 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  _T_1782_1 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  _T_1783_0 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  _T_1783_1 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  _T_1794_0 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  _T_1794_1 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  _T_1795_0 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  _T_1795_1 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  _T_1806_0 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  _T_1806_1 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  _T_1807_0 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  _T_1807_1 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  _T_1818_0 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  _T_1818_1 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  _T_1819_0 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  _T_1819_1 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  _T_1831_0 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  _T_1831_1 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  _T_1843_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  _T_1843_1 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  _T_1855_0 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  _T_1855_1 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  _T_1866_0 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  _T_1866_1 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  _T_1867_0 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  _T_1867_1 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  _T_1878_0 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  _T_1878_1 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  _T_1879_0 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  _T_1879_1 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  _T_1890_0 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  _T_1890_1 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  _T_1891_0 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  _T_1891_1 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  _T_1903_0 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  _T_1903_1 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  _T_1915_0 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  _T_1915_1 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  _T_1927_0 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  _T_1927_1 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  _T_1939_0 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  _T_1939_1 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  _T_1951_0 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  _T_1951_1 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  _T_1963_0 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  _T_1963_1 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  _T_1975_0 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  _T_1975_1 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  _T_1987_0 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  _T_1987_1 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  _T_1999_0 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  _T_1999_1 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  _T_2011_0 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  _T_2011_1 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  _T_2023_0 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  _T_2023_1 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  _T_2035_0 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  _T_2035_1 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  _T_2047_0 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  _T_2047_1 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  _T_2059_0 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  _T_2059_1 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  _T_2071_0 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  _T_2071_1 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  _T_2083_0 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  _T_2083_1 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  _T_2095_0 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  _T_2095_1 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  _T_2107_0 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  _T_2107_1 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  _T_2119_0 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  _T_2119_1 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  _T_2131_0 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  _T_2131_1 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  _T_2143_0 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  _T_2143_1 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  _T_2155_0 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  _T_2155_1 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  _T_2167_0 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  _T_2167_1 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  _T_2179_0 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  _T_2179_1 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  _T_2191_0 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  _T_2191_1 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  _T_2203_0 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  _T_2203_1 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  _T_2215_0 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  _T_2215_1 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  _T_2227_0 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  _T_2227_1 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  _T_2239_0 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  _T_2239_1 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  _T_2251_0 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  _T_2251_1 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  _T_2263_0 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  _T_2263_1 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  _T_2275_0 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  _T_2275_1 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  _T_2287_0 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  _T_2287_1 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  _T_2299_0 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  _T_2299_1 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  _T_2311_0 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  _T_2311_1 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  _T_2323_0 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  _T_2323_1 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  _T_2335_0 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  _T_2335_1 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  _T_2347_0 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  _T_2347_1 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  _T_2359_0 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  _T_2359_1 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  _T_2371_0 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  _T_2371_1 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  _T_2383_0 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  _T_2383_1 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  _T_2395_0 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  _T_2395_1 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  _T_2407_0 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  _T_2407_1 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  _T_2419_0 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  _T_2419_1 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  _T_2431_0 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  _T_2431_1 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  _T_2443_0 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  _T_2443_1 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  _T_2455_0 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  _T_2455_1 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  _T_2467_0 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  _T_2467_1 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  _T_2479_0 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  _T_2479_1 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  _T_2491_0 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  _T_2491_1 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  _T_2503_0 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  _T_2503_1 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  _T_2515_0 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  _T_2515_1 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  _T_2527_0 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  _T_2527_1 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  _T_2539_0 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  _T_2539_1 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  _T_2551_0 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  _T_2551_1 = _RAND_741[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= io_pixelColorBack;
    pixelColorBackReg <= _T;
    _T_3_0 <= _T_3_1;
    _T_3_1 <= io_spriteVisibleReg_0;
    _T_4_0 <= _T_4_1;
    _T_4_1 <= io_inSprite_0;
    _T_11_0 <= _T_11_1;
    _T_11_1 <= io_spriteVisibleReg_1;
    _T_12_0 <= _T_12_1;
    _T_12_1 <= io_inSprite_1;
    _T_19_0 <= _T_19_1;
    _T_19_1 <= io_spriteVisibleReg_2;
    _T_20_0 <= _T_20_1;
    _T_20_1 <= io_inSprite_2;
    _T_27_0 <= _T_27_1;
    _T_27_1 <= io_spriteVisibleReg_3;
    _T_28_0 <= _T_28_1;
    _T_28_1 <= io_inSprite_3;
    _T_35_0 <= _T_35_1;
    _T_35_1 <= io_spriteVisibleReg_4;
    _T_36_0 <= _T_36_1;
    _T_36_1 <= io_inSprite_4;
    _T_43_0 <= _T_43_1;
    _T_43_1 <= io_spriteVisibleReg_5;
    _T_44_0 <= _T_44_1;
    _T_44_1 <= io_inSprite_5;
    _T_51_0 <= _T_51_1;
    _T_51_1 <= io_spriteVisibleReg_6;
    _T_52_0 <= _T_52_1;
    _T_52_1 <= io_inSprite_6;
    _T_59_0 <= _T_59_1;
    _T_59_1 <= io_spriteVisibleReg_7;
    _T_60_0 <= _T_60_1;
    _T_60_1 <= io_inSprite_7;
    _T_67_0 <= _T_67_1;
    _T_67_1 <= io_spriteVisibleReg_8;
    _T_68_0 <= _T_68_1;
    _T_68_1 <= io_inSprite_8;
    _T_75_0 <= _T_75_1;
    _T_75_1 <= io_spriteVisibleReg_9;
    _T_76_0 <= _T_76_1;
    _T_76_1 <= io_inSprite_9;
    _T_83_0 <= _T_83_1;
    _T_83_1 <= io_spriteVisibleReg_10;
    _T_84_0 <= _T_84_1;
    _T_84_1 <= io_inSprite_10;
    _T_91_0 <= _T_91_1;
    _T_91_1 <= io_spriteVisibleReg_11;
    _T_92_0 <= _T_92_1;
    _T_92_1 <= io_inSprite_11;
    _T_99_0 <= _T_99_1;
    _T_99_1 <= io_spriteVisibleReg_12;
    _T_100_0 <= _T_100_1;
    _T_100_1 <= io_inSprite_12;
    _T_107_0 <= _T_107_1;
    _T_107_1 <= io_spriteVisibleReg_13;
    _T_108_0 <= _T_108_1;
    _T_108_1 <= io_inSprite_13;
    _T_115_0 <= _T_115_1;
    _T_115_1 <= io_spriteVisibleReg_14;
    _T_116_0 <= _T_116_1;
    _T_116_1 <= io_inSprite_14;
    _T_123_0 <= _T_123_1;
    _T_123_1 <= io_spriteVisibleReg_15;
    _T_124_0 <= _T_124_1;
    _T_124_1 <= io_inSprite_15;
    _T_131_0 <= _T_131_1;
    _T_131_1 <= io_spriteVisibleReg_16;
    _T_132_0 <= _T_132_1;
    _T_132_1 <= io_inSprite_16;
    _T_139_0 <= _T_139_1;
    _T_139_1 <= io_spriteVisibleReg_17;
    _T_140_0 <= _T_140_1;
    _T_140_1 <= io_inSprite_17;
    _T_147_0 <= _T_147_1;
    _T_147_1 <= io_spriteVisibleReg_18;
    _T_148_0 <= _T_148_1;
    _T_148_1 <= io_inSprite_18;
    _T_155_0 <= _T_155_1;
    _T_155_1 <= io_spriteVisibleReg_19;
    _T_156_0 <= _T_156_1;
    _T_156_1 <= io_inSprite_19;
    _T_163_0 <= _T_163_1;
    _T_163_1 <= io_spriteVisibleReg_20;
    _T_164_0 <= _T_164_1;
    _T_164_1 <= io_inSprite_20;
    _T_171_0 <= _T_171_1;
    _T_171_1 <= io_spriteVisibleReg_21;
    _T_172_0 <= _T_172_1;
    _T_172_1 <= io_inSprite_21;
    _T_179_0 <= _T_179_1;
    _T_179_1 <= io_spriteVisibleReg_22;
    _T_180_0 <= _T_180_1;
    _T_180_1 <= io_inSprite_22;
    _T_187_0 <= _T_187_1;
    _T_187_1 <= io_spriteVisibleReg_23;
    _T_188_0 <= _T_188_1;
    _T_188_1 <= io_inSprite_23;
    _T_195_0 <= _T_195_1;
    _T_195_1 <= io_spriteVisibleReg_24;
    _T_196_0 <= _T_196_1;
    _T_196_1 <= io_inSprite_24;
    _T_203_0 <= _T_203_1;
    _T_203_1 <= io_spriteVisibleReg_25;
    _T_204_0 <= _T_204_1;
    _T_204_1 <= io_inSprite_25;
    _T_211_0 <= _T_211_1;
    _T_211_1 <= io_spriteVisibleReg_26;
    _T_212_0 <= _T_212_1;
    _T_212_1 <= io_inSprite_26;
    _T_219_0 <= _T_219_1;
    _T_219_1 <= io_spriteVisibleReg_27;
    _T_220_0 <= _T_220_1;
    _T_220_1 <= io_inSprite_27;
    _T_227_0 <= _T_227_1;
    _T_227_1 <= io_spriteVisibleReg_28;
    _T_228_0 <= _T_228_1;
    _T_228_1 <= io_inSprite_28;
    _T_235_0 <= _T_235_1;
    _T_235_1 <= io_spriteVisibleReg_29;
    _T_236_0 <= _T_236_1;
    _T_236_1 <= io_inSprite_29;
    _T_243_0 <= _T_243_1;
    _T_243_1 <= io_spriteVisibleReg_30;
    _T_244_0 <= _T_244_1;
    _T_244_1 <= io_inSprite_30;
    _T_251_0 <= _T_251_1;
    _T_251_1 <= io_spriteVisibleReg_31;
    _T_252_0 <= _T_252_1;
    _T_252_1 <= io_inSprite_31;
    _T_259_0 <= _T_259_1;
    _T_259_1 <= io_spriteVisibleReg_32;
    _T_260_0 <= _T_260_1;
    _T_260_1 <= io_inSprite_32;
    _T_267_0 <= _T_267_1;
    _T_267_1 <= io_spriteVisibleReg_33;
    _T_268_0 <= _T_268_1;
    _T_268_1 <= io_inSprite_33;
    _T_276_0 <= _T_276_1;
    _T_276_1 <= io_inSprite_34;
    _T_284_0 <= _T_284_1;
    _T_284_1 <= io_inSprite_35;
    _T_292_0 <= _T_292_1;
    _T_292_1 <= io_inSprite_36;
    _T_300_0 <= _T_300_1;
    _T_300_1 <= io_inSprite_37;
    _T_308_0 <= _T_308_1;
    _T_308_1 <= io_inSprite_38;
    _T_316_0 <= _T_316_1;
    _T_316_1 <= io_inSprite_39;
    _T_324_0 <= _T_324_1;
    _T_324_1 <= io_inSprite_40;
    _T_331_0 <= _T_331_1;
    _T_331_1 <= io_spriteVisibleReg_41;
    _T_332_0 <= _T_332_1;
    _T_332_1 <= io_inSprite_41;
    _T_339_0 <= _T_339_1;
    _T_339_1 <= io_spriteVisibleReg_42;
    _T_340_0 <= _T_340_1;
    _T_340_1 <= io_inSprite_42;
    _T_347_0 <= _T_347_1;
    _T_347_1 <= io_spriteVisibleReg_43;
    _T_348_0 <= _T_348_1;
    _T_348_1 <= io_inSprite_43;
    _T_355_0 <= _T_355_1;
    _T_355_1 <= io_spriteVisibleReg_44;
    _T_356_0 <= _T_356_1;
    _T_356_1 <= io_inSprite_44;
    _T_363_0 <= _T_363_1;
    _T_363_1 <= io_spriteVisibleReg_45;
    _T_364_0 <= _T_364_1;
    _T_364_1 <= io_inSprite_45;
    _T_371_0 <= _T_371_1;
    _T_371_1 <= io_spriteVisibleReg_46;
    _T_372_0 <= _T_372_1;
    _T_372_1 <= io_inSprite_46;
    _T_379_0 <= _T_379_1;
    _T_379_1 <= io_spriteVisibleReg_47;
    _T_380_0 <= _T_380_1;
    _T_380_1 <= io_inSprite_47;
    _T_387_0 <= _T_387_1;
    _T_387_1 <= io_spriteVisibleReg_48;
    _T_388_0 <= _T_388_1;
    _T_388_1 <= io_inSprite_48;
    _T_395_0 <= _T_395_1;
    _T_395_1 <= io_spriteVisibleReg_49;
    _T_396_0 <= _T_396_1;
    _T_396_1 <= io_inSprite_49;
    _T_403_0 <= _T_403_1;
    _T_403_1 <= io_spriteVisibleReg_50;
    _T_404_0 <= _T_404_1;
    _T_404_1 <= io_inSprite_50;
    _T_411_0 <= _T_411_1;
    _T_411_1 <= io_spriteVisibleReg_51;
    _T_412_0 <= _T_412_1;
    _T_412_1 <= io_inSprite_51;
    _T_420_0 <= _T_420_1;
    _T_420_1 <= io_inSprite_52;
    _T_428_0 <= _T_428_1;
    _T_428_1 <= io_inSprite_53;
    _T_436_0 <= _T_436_1;
    _T_436_1 <= io_inSprite_54;
    _T_443_0 <= _T_443_1;
    _T_443_1 <= io_spriteVisibleReg_55;
    _T_444_0 <= _T_444_1;
    _T_444_1 <= io_inSprite_55;
    _T_451_0 <= _T_451_1;
    _T_451_1 <= io_spriteVisibleReg_56;
    _T_452_0 <= _T_452_1;
    _T_452_1 <= io_inSprite_56;
    _T_459_0 <= _T_459_1;
    _T_459_1 <= io_spriteVisibleReg_57;
    _T_460_0 <= _T_460_1;
    _T_460_1 <= io_inSprite_57;
    _T_468_0 <= _T_468_1;
    _T_468_1 <= io_inSprite_58;
    _T_476_0 <= _T_476_1;
    _T_476_1 <= io_inSprite_59;
    _T_484_0 <= _T_484_1;
    _T_484_1 <= io_inSprite_60;
    _T_491_0 <= _T_491_1;
    _T_491_1 <= io_spriteVisibleReg_61;
    _T_492_0 <= _T_492_1;
    _T_492_1 <= io_inSprite_61;
    _T_499_0 <= _T_499_1;
    _T_499_1 <= io_spriteVisibleReg_62;
    _T_500_0 <= _T_500_1;
    _T_500_1 <= io_inSprite_62;
    _T_507_0 <= _T_507_1;
    _T_507_1 <= io_spriteVisibleReg_63;
    _T_508_0 <= _T_508_1;
    _T_508_1 <= io_inSprite_63;
    _T_515_0 <= _T_515_1;
    _T_515_1 <= io_spriteVisibleReg_64;
    _T_516_0 <= _T_516_1;
    _T_516_1 <= io_inSprite_64;
    _T_523_0 <= _T_523_1;
    _T_523_1 <= io_spriteVisibleReg_65;
    _T_524_0 <= _T_524_1;
    _T_524_1 <= io_inSprite_65;
    _T_531_0 <= _T_531_1;
    _T_531_1 <= io_spriteVisibleReg_66;
    _T_532_0 <= _T_532_1;
    _T_532_1 <= io_inSprite_66;
    _T_540_0 <= _T_540_1;
    _T_540_1 <= io_inSprite_67;
    _T_548_0 <= _T_548_1;
    _T_548_1 <= io_inSprite_68;
    _T_556_0 <= _T_556_1;
    _T_556_1 <= io_inSprite_69;
    _T_563_0 <= _T_563_1;
    _T_563_1 <= io_spriteVisibleReg_70;
    _T_564_0 <= _T_564_1;
    _T_564_1 <= io_inSprite_70;
    _T_571_0 <= _T_571_1;
    _T_571_1 <= io_spriteVisibleReg_71;
    _T_572_0 <= _T_572_1;
    _T_572_1 <= io_inSprite_71;
    _T_579_0 <= _T_579_1;
    _T_579_1 <= io_spriteVisibleReg_72;
    _T_580_0 <= _T_580_1;
    _T_580_1 <= io_inSprite_72;
    _T_588_0 <= _T_588_1;
    _T_588_1 <= io_inSprite_73;
    _T_596_0 <= _T_596_1;
    _T_596_1 <= io_inSprite_74;
    _T_604_0 <= _T_604_1;
    _T_604_1 <= io_inSprite_75;
    _T_612_0 <= _T_612_1;
    _T_612_1 <= io_inSprite_76;
    _T_620_0 <= _T_620_1;
    _T_620_1 <= io_inSprite_77;
    _T_628_0 <= _T_628_1;
    _T_628_1 <= io_inSprite_78;
    _T_636_0 <= _T_636_1;
    _T_636_1 <= io_inSprite_79;
    _T_644_0 <= _T_644_1;
    _T_644_1 <= io_inSprite_80;
    _T_652_0 <= _T_652_1;
    _T_652_1 <= io_inSprite_81;
    _T_660_0 <= _T_660_1;
    _T_660_1 <= io_inSprite_82;
    _T_668_0 <= _T_668_1;
    _T_668_1 <= io_inSprite_83;
    _T_676_0 <= _T_676_1;
    _T_676_1 <= io_inSprite_84;
    _T_684_0 <= _T_684_1;
    _T_684_1 <= io_inSprite_85;
    _T_692_0 <= _T_692_1;
    _T_692_1 <= io_inSprite_86;
    _T_700_0 <= _T_700_1;
    _T_700_1 <= io_inSprite_87;
    _T_708_0 <= _T_708_1;
    _T_708_1 <= io_inSprite_88;
    _T_716_0 <= _T_716_1;
    _T_716_1 <= io_inSprite_89;
    _T_724_0 <= _T_724_1;
    _T_724_1 <= io_inSprite_90;
    _T_732_0 <= _T_732_1;
    _T_732_1 <= io_inSprite_91;
    _T_740_0 <= _T_740_1;
    _T_740_1 <= io_inSprite_92;
    _T_748_0 <= _T_748_1;
    _T_748_1 <= io_inSprite_93;
    _T_756_0 <= _T_756_1;
    _T_756_1 <= io_inSprite_94;
    _T_764_0 <= _T_764_1;
    _T_764_1 <= io_inSprite_95;
    _T_772_0 <= _T_772_1;
    _T_772_1 <= io_inSprite_96;
    _T_780_0 <= _T_780_1;
    _T_780_1 <= io_inSprite_97;
    _T_788_0 <= _T_788_1;
    _T_788_1 <= io_inSprite_98;
    _T_796_0 <= _T_796_1;
    _T_796_1 <= io_inSprite_99;
    _T_804_0 <= _T_804_1;
    _T_804_1 <= io_inSprite_100;
    _T_812_0 <= _T_812_1;
    _T_812_1 <= io_inSprite_101;
    _T_820_0 <= _T_820_1;
    _T_820_1 <= io_inSprite_102;
    _T_828_0 <= _T_828_1;
    _T_828_1 <= io_inSprite_103;
    _T_836_0 <= _T_836_1;
    _T_836_1 <= io_inSprite_104;
    _T_844_0 <= _T_844_1;
    _T_844_1 <= io_inSprite_105;
    _T_852_0 <= _T_852_1;
    _T_852_1 <= io_inSprite_106;
    _T_860_0 <= _T_860_1;
    _T_860_1 <= io_inSprite_107;
    _T_868_0 <= _T_868_1;
    _T_868_1 <= io_inSprite_108;
    _T_876_0 <= _T_876_1;
    _T_876_1 <= io_inSprite_109;
    _T_884_0 <= _T_884_1;
    _T_884_1 <= io_inSprite_110;
    _T_892_0 <= _T_892_1;
    _T_892_1 <= io_inSprite_111;
    _T_900_0 <= _T_900_1;
    _T_900_1 <= io_inSprite_112;
    _T_908_0 <= _T_908_1;
    _T_908_1 <= io_inSprite_113;
    _T_916_0 <= _T_916_1;
    _T_916_1 <= io_inSprite_114;
    _T_924_0 <= _T_924_1;
    _T_924_1 <= io_inSprite_115;
    _T_932_0 <= _T_932_1;
    _T_932_1 <= io_inSprite_116;
    _T_940_0 <= _T_940_1;
    _T_940_1 <= io_inSprite_117;
    _T_948_0 <= _T_948_1;
    _T_948_1 <= io_inSprite_118;
    _T_956_0 <= _T_956_1;
    _T_956_1 <= io_inSprite_119;
    _T_964_0 <= _T_964_1;
    _T_964_1 <= io_inSprite_120;
    _T_972_0 <= _T_972_1;
    _T_972_1 <= io_inSprite_121;
    _T_980_0 <= _T_980_1;
    _T_980_1 <= io_inSprite_122;
    _T_988_0 <= _T_988_1;
    _T_988_1 <= io_inSprite_123;
    _T_996_0 <= _T_996_1;
    _T_996_1 <= io_inSprite_124;
    _T_1004_0 <= _T_1004_1;
    _T_1004_1 <= io_inSprite_125;
    _T_1012_0 <= _T_1012_1;
    _T_1012_1 <= io_inSprite_126;
    _T_1020_0 <= _T_1020_1;
    _T_1020_1 <= io_inSprite_127;
    _T_1026_0 <= _T_1026_1;
    _T_1026_1 <= io_spriteVisibleReg_0;
    _T_1027_0 <= _T_1027_1;
    _T_1027_1 <= io_inSprite_0;
    _T_1038_0 <= _T_1038_1;
    _T_1038_1 <= io_spriteVisibleReg_1;
    _T_1039_0 <= _T_1039_1;
    _T_1039_1 <= io_inSprite_1;
    _T_1050_0 <= _T_1050_1;
    _T_1050_1 <= io_spriteVisibleReg_2;
    _T_1051_0 <= _T_1051_1;
    _T_1051_1 <= io_inSprite_2;
    _T_1062_0 <= _T_1062_1;
    _T_1062_1 <= io_spriteVisibleReg_3;
    _T_1063_0 <= _T_1063_1;
    _T_1063_1 <= io_inSprite_3;
    _T_1074_0 <= _T_1074_1;
    _T_1074_1 <= io_spriteVisibleReg_4;
    _T_1075_0 <= _T_1075_1;
    _T_1075_1 <= io_inSprite_4;
    _T_1086_0 <= _T_1086_1;
    _T_1086_1 <= io_spriteVisibleReg_5;
    _T_1087_0 <= _T_1087_1;
    _T_1087_1 <= io_inSprite_5;
    _T_1098_0 <= _T_1098_1;
    _T_1098_1 <= io_spriteVisibleReg_6;
    _T_1099_0 <= _T_1099_1;
    _T_1099_1 <= io_inSprite_6;
    _T_1110_0 <= _T_1110_1;
    _T_1110_1 <= io_spriteVisibleReg_7;
    _T_1111_0 <= _T_1111_1;
    _T_1111_1 <= io_inSprite_7;
    _T_1122_0 <= _T_1122_1;
    _T_1122_1 <= io_spriteVisibleReg_8;
    _T_1123_0 <= _T_1123_1;
    _T_1123_1 <= io_inSprite_8;
    _T_1134_0 <= _T_1134_1;
    _T_1134_1 <= io_spriteVisibleReg_9;
    _T_1135_0 <= _T_1135_1;
    _T_1135_1 <= io_inSprite_9;
    _T_1146_0 <= _T_1146_1;
    _T_1146_1 <= io_spriteVisibleReg_10;
    _T_1147_0 <= _T_1147_1;
    _T_1147_1 <= io_inSprite_10;
    _T_1158_0 <= _T_1158_1;
    _T_1158_1 <= io_spriteVisibleReg_11;
    _T_1159_0 <= _T_1159_1;
    _T_1159_1 <= io_inSprite_11;
    _T_1170_0 <= _T_1170_1;
    _T_1170_1 <= io_spriteVisibleReg_12;
    _T_1171_0 <= _T_1171_1;
    _T_1171_1 <= io_inSprite_12;
    _T_1182_0 <= _T_1182_1;
    _T_1182_1 <= io_spriteVisibleReg_13;
    _T_1183_0 <= _T_1183_1;
    _T_1183_1 <= io_inSprite_13;
    _T_1194_0 <= _T_1194_1;
    _T_1194_1 <= io_spriteVisibleReg_14;
    _T_1195_0 <= _T_1195_1;
    _T_1195_1 <= io_inSprite_14;
    _T_1206_0 <= _T_1206_1;
    _T_1206_1 <= io_spriteVisibleReg_15;
    _T_1207_0 <= _T_1207_1;
    _T_1207_1 <= io_inSprite_15;
    _T_1218_0 <= _T_1218_1;
    _T_1218_1 <= io_spriteVisibleReg_16;
    _T_1219_0 <= _T_1219_1;
    _T_1219_1 <= io_inSprite_16;
    _T_1230_0 <= _T_1230_1;
    _T_1230_1 <= io_spriteVisibleReg_17;
    _T_1231_0 <= _T_1231_1;
    _T_1231_1 <= io_inSprite_17;
    _T_1242_0 <= _T_1242_1;
    _T_1242_1 <= io_spriteVisibleReg_18;
    _T_1243_0 <= _T_1243_1;
    _T_1243_1 <= io_inSprite_18;
    _T_1254_0 <= _T_1254_1;
    _T_1254_1 <= io_spriteVisibleReg_19;
    _T_1255_0 <= _T_1255_1;
    _T_1255_1 <= io_inSprite_19;
    _T_1266_0 <= _T_1266_1;
    _T_1266_1 <= io_spriteVisibleReg_20;
    _T_1267_0 <= _T_1267_1;
    _T_1267_1 <= io_inSprite_20;
    _T_1278_0 <= _T_1278_1;
    _T_1278_1 <= io_spriteVisibleReg_21;
    _T_1279_0 <= _T_1279_1;
    _T_1279_1 <= io_inSprite_21;
    _T_1290_0 <= _T_1290_1;
    _T_1290_1 <= io_spriteVisibleReg_22;
    _T_1291_0 <= _T_1291_1;
    _T_1291_1 <= io_inSprite_22;
    _T_1302_0 <= _T_1302_1;
    _T_1302_1 <= io_spriteVisibleReg_23;
    _T_1303_0 <= _T_1303_1;
    _T_1303_1 <= io_inSprite_23;
    _T_1314_0 <= _T_1314_1;
    _T_1314_1 <= io_spriteVisibleReg_24;
    _T_1315_0 <= _T_1315_1;
    _T_1315_1 <= io_inSprite_24;
    _T_1326_0 <= _T_1326_1;
    _T_1326_1 <= io_spriteVisibleReg_25;
    _T_1327_0 <= _T_1327_1;
    _T_1327_1 <= io_inSprite_25;
    _T_1338_0 <= _T_1338_1;
    _T_1338_1 <= io_spriteVisibleReg_26;
    _T_1339_0 <= _T_1339_1;
    _T_1339_1 <= io_inSprite_26;
    _T_1350_0 <= _T_1350_1;
    _T_1350_1 <= io_spriteVisibleReg_27;
    _T_1351_0 <= _T_1351_1;
    _T_1351_1 <= io_inSprite_27;
    _T_1362_0 <= _T_1362_1;
    _T_1362_1 <= io_spriteVisibleReg_28;
    _T_1363_0 <= _T_1363_1;
    _T_1363_1 <= io_inSprite_28;
    _T_1374_0 <= _T_1374_1;
    _T_1374_1 <= io_spriteVisibleReg_29;
    _T_1375_0 <= _T_1375_1;
    _T_1375_1 <= io_inSprite_29;
    _T_1386_0 <= _T_1386_1;
    _T_1386_1 <= io_spriteVisibleReg_30;
    _T_1387_0 <= _T_1387_1;
    _T_1387_1 <= io_inSprite_30;
    _T_1398_0 <= _T_1398_1;
    _T_1398_1 <= io_spriteVisibleReg_31;
    _T_1399_0 <= _T_1399_1;
    _T_1399_1 <= io_inSprite_31;
    _T_1410_0 <= _T_1410_1;
    _T_1410_1 <= io_spriteVisibleReg_32;
    _T_1411_0 <= _T_1411_1;
    _T_1411_1 <= io_inSprite_32;
    _T_1422_0 <= _T_1422_1;
    _T_1422_1 <= io_spriteVisibleReg_33;
    _T_1423_0 <= _T_1423_1;
    _T_1423_1 <= io_inSprite_33;
    _T_1435_0 <= _T_1435_1;
    _T_1435_1 <= io_inSprite_34;
    _T_1447_0 <= _T_1447_1;
    _T_1447_1 <= io_inSprite_35;
    _T_1459_0 <= _T_1459_1;
    _T_1459_1 <= io_inSprite_36;
    _T_1471_0 <= _T_1471_1;
    _T_1471_1 <= io_inSprite_37;
    _T_1483_0 <= _T_1483_1;
    _T_1483_1 <= io_inSprite_38;
    _T_1495_0 <= _T_1495_1;
    _T_1495_1 <= io_inSprite_39;
    _T_1507_0 <= _T_1507_1;
    _T_1507_1 <= io_inSprite_40;
    _T_1518_0 <= _T_1518_1;
    _T_1518_1 <= io_spriteVisibleReg_41;
    _T_1519_0 <= _T_1519_1;
    _T_1519_1 <= io_inSprite_41;
    _T_1530_0 <= _T_1530_1;
    _T_1530_1 <= io_spriteVisibleReg_42;
    _T_1531_0 <= _T_1531_1;
    _T_1531_1 <= io_inSprite_42;
    _T_1542_0 <= _T_1542_1;
    _T_1542_1 <= io_spriteVisibleReg_43;
    _T_1543_0 <= _T_1543_1;
    _T_1543_1 <= io_inSprite_43;
    _T_1554_0 <= _T_1554_1;
    _T_1554_1 <= io_spriteVisibleReg_44;
    _T_1555_0 <= _T_1555_1;
    _T_1555_1 <= io_inSprite_44;
    _T_1566_0 <= _T_1566_1;
    _T_1566_1 <= io_spriteVisibleReg_45;
    _T_1567_0 <= _T_1567_1;
    _T_1567_1 <= io_inSprite_45;
    _T_1578_0 <= _T_1578_1;
    _T_1578_1 <= io_spriteVisibleReg_46;
    _T_1579_0 <= _T_1579_1;
    _T_1579_1 <= io_inSprite_46;
    _T_1590_0 <= _T_1590_1;
    _T_1590_1 <= io_spriteVisibleReg_47;
    _T_1591_0 <= _T_1591_1;
    _T_1591_1 <= io_inSprite_47;
    _T_1602_0 <= _T_1602_1;
    _T_1602_1 <= io_spriteVisibleReg_48;
    _T_1603_0 <= _T_1603_1;
    _T_1603_1 <= io_inSprite_48;
    _T_1614_0 <= _T_1614_1;
    _T_1614_1 <= io_spriteVisibleReg_49;
    _T_1615_0 <= _T_1615_1;
    _T_1615_1 <= io_inSprite_49;
    _T_1626_0 <= _T_1626_1;
    _T_1626_1 <= io_spriteVisibleReg_50;
    _T_1627_0 <= _T_1627_1;
    _T_1627_1 <= io_inSprite_50;
    _T_1638_0 <= _T_1638_1;
    _T_1638_1 <= io_spriteVisibleReg_51;
    _T_1639_0 <= _T_1639_1;
    _T_1639_1 <= io_inSprite_51;
    _T_1651_0 <= _T_1651_1;
    _T_1651_1 <= io_inSprite_52;
    _T_1663_0 <= _T_1663_1;
    _T_1663_1 <= io_inSprite_53;
    _T_1675_0 <= _T_1675_1;
    _T_1675_1 <= io_inSprite_54;
    _T_1686_0 <= _T_1686_1;
    _T_1686_1 <= io_spriteVisibleReg_55;
    _T_1687_0 <= _T_1687_1;
    _T_1687_1 <= io_inSprite_55;
    _T_1698_0 <= _T_1698_1;
    _T_1698_1 <= io_spriteVisibleReg_56;
    _T_1699_0 <= _T_1699_1;
    _T_1699_1 <= io_inSprite_56;
    _T_1710_0 <= _T_1710_1;
    _T_1710_1 <= io_spriteVisibleReg_57;
    _T_1711_0 <= _T_1711_1;
    _T_1711_1 <= io_inSprite_57;
    _T_1723_0 <= _T_1723_1;
    _T_1723_1 <= io_inSprite_58;
    _T_1735_0 <= _T_1735_1;
    _T_1735_1 <= io_inSprite_59;
    _T_1747_0 <= _T_1747_1;
    _T_1747_1 <= io_inSprite_60;
    _T_1758_0 <= _T_1758_1;
    _T_1758_1 <= io_spriteVisibleReg_61;
    _T_1759_0 <= _T_1759_1;
    _T_1759_1 <= io_inSprite_61;
    _T_1770_0 <= _T_1770_1;
    _T_1770_1 <= io_spriteVisibleReg_62;
    _T_1771_0 <= _T_1771_1;
    _T_1771_1 <= io_inSprite_62;
    _T_1782_0 <= _T_1782_1;
    _T_1782_1 <= io_spriteVisibleReg_63;
    _T_1783_0 <= _T_1783_1;
    _T_1783_1 <= io_inSprite_63;
    _T_1794_0 <= _T_1794_1;
    _T_1794_1 <= io_spriteVisibleReg_64;
    _T_1795_0 <= _T_1795_1;
    _T_1795_1 <= io_inSprite_64;
    _T_1806_0 <= _T_1806_1;
    _T_1806_1 <= io_spriteVisibleReg_65;
    _T_1807_0 <= _T_1807_1;
    _T_1807_1 <= io_inSprite_65;
    _T_1818_0 <= _T_1818_1;
    _T_1818_1 <= io_spriteVisibleReg_66;
    _T_1819_0 <= _T_1819_1;
    _T_1819_1 <= io_inSprite_66;
    _T_1831_0 <= _T_1831_1;
    _T_1831_1 <= io_inSprite_67;
    _T_1843_0 <= _T_1843_1;
    _T_1843_1 <= io_inSprite_68;
    _T_1855_0 <= _T_1855_1;
    _T_1855_1 <= io_inSprite_69;
    _T_1866_0 <= _T_1866_1;
    _T_1866_1 <= io_spriteVisibleReg_70;
    _T_1867_0 <= _T_1867_1;
    _T_1867_1 <= io_inSprite_70;
    _T_1878_0 <= _T_1878_1;
    _T_1878_1 <= io_spriteVisibleReg_71;
    _T_1879_0 <= _T_1879_1;
    _T_1879_1 <= io_inSprite_71;
    _T_1890_0 <= _T_1890_1;
    _T_1890_1 <= io_spriteVisibleReg_72;
    _T_1891_0 <= _T_1891_1;
    _T_1891_1 <= io_inSprite_72;
    _T_1903_0 <= _T_1903_1;
    _T_1903_1 <= io_inSprite_73;
    _T_1915_0 <= _T_1915_1;
    _T_1915_1 <= io_inSprite_74;
    _T_1927_0 <= _T_1927_1;
    _T_1927_1 <= io_inSprite_75;
    _T_1939_0 <= _T_1939_1;
    _T_1939_1 <= io_inSprite_76;
    _T_1951_0 <= _T_1951_1;
    _T_1951_1 <= io_inSprite_77;
    _T_1963_0 <= _T_1963_1;
    _T_1963_1 <= io_inSprite_78;
    _T_1975_0 <= _T_1975_1;
    _T_1975_1 <= io_inSprite_79;
    _T_1987_0 <= _T_1987_1;
    _T_1987_1 <= io_inSprite_80;
    _T_1999_0 <= _T_1999_1;
    _T_1999_1 <= io_inSprite_81;
    _T_2011_0 <= _T_2011_1;
    _T_2011_1 <= io_inSprite_82;
    _T_2023_0 <= _T_2023_1;
    _T_2023_1 <= io_inSprite_83;
    _T_2035_0 <= _T_2035_1;
    _T_2035_1 <= io_inSprite_84;
    _T_2047_0 <= _T_2047_1;
    _T_2047_1 <= io_inSprite_85;
    _T_2059_0 <= _T_2059_1;
    _T_2059_1 <= io_inSprite_86;
    _T_2071_0 <= _T_2071_1;
    _T_2071_1 <= io_inSprite_87;
    _T_2083_0 <= _T_2083_1;
    _T_2083_1 <= io_inSprite_88;
    _T_2095_0 <= _T_2095_1;
    _T_2095_1 <= io_inSprite_89;
    _T_2107_0 <= _T_2107_1;
    _T_2107_1 <= io_inSprite_90;
    _T_2119_0 <= _T_2119_1;
    _T_2119_1 <= io_inSprite_91;
    _T_2131_0 <= _T_2131_1;
    _T_2131_1 <= io_inSprite_92;
    _T_2143_0 <= _T_2143_1;
    _T_2143_1 <= io_inSprite_93;
    _T_2155_0 <= _T_2155_1;
    _T_2155_1 <= io_inSprite_94;
    _T_2167_0 <= _T_2167_1;
    _T_2167_1 <= io_inSprite_95;
    _T_2179_0 <= _T_2179_1;
    _T_2179_1 <= io_inSprite_96;
    _T_2191_0 <= _T_2191_1;
    _T_2191_1 <= io_inSprite_97;
    _T_2203_0 <= _T_2203_1;
    _T_2203_1 <= io_inSprite_98;
    _T_2215_0 <= _T_2215_1;
    _T_2215_1 <= io_inSprite_99;
    _T_2227_0 <= _T_2227_1;
    _T_2227_1 <= io_inSprite_100;
    _T_2239_0 <= _T_2239_1;
    _T_2239_1 <= io_inSprite_101;
    _T_2251_0 <= _T_2251_1;
    _T_2251_1 <= io_inSprite_102;
    _T_2263_0 <= _T_2263_1;
    _T_2263_1 <= io_inSprite_103;
    _T_2275_0 <= _T_2275_1;
    _T_2275_1 <= io_inSprite_104;
    _T_2287_0 <= _T_2287_1;
    _T_2287_1 <= io_inSprite_105;
    _T_2299_0 <= _T_2299_1;
    _T_2299_1 <= io_inSprite_106;
    _T_2311_0 <= _T_2311_1;
    _T_2311_1 <= io_inSprite_107;
    _T_2323_0 <= _T_2323_1;
    _T_2323_1 <= io_inSprite_108;
    _T_2335_0 <= _T_2335_1;
    _T_2335_1 <= io_inSprite_109;
    _T_2347_0 <= _T_2347_1;
    _T_2347_1 <= io_inSprite_110;
    _T_2359_0 <= _T_2359_1;
    _T_2359_1 <= io_inSprite_111;
    _T_2371_0 <= _T_2371_1;
    _T_2371_1 <= io_inSprite_112;
    _T_2383_0 <= _T_2383_1;
    _T_2383_1 <= io_inSprite_113;
    _T_2395_0 <= _T_2395_1;
    _T_2395_1 <= io_inSprite_114;
    _T_2407_0 <= _T_2407_1;
    _T_2407_1 <= io_inSprite_115;
    _T_2419_0 <= _T_2419_1;
    _T_2419_1 <= io_inSprite_116;
    _T_2431_0 <= _T_2431_1;
    _T_2431_1 <= io_inSprite_117;
    _T_2443_0 <= _T_2443_1;
    _T_2443_1 <= io_inSprite_118;
    _T_2455_0 <= _T_2455_1;
    _T_2455_1 <= io_inSprite_119;
    _T_2467_0 <= _T_2467_1;
    _T_2467_1 <= io_inSprite_120;
    _T_2479_0 <= _T_2479_1;
    _T_2479_1 <= io_inSprite_121;
    _T_2491_0 <= _T_2491_1;
    _T_2491_1 <= io_inSprite_122;
    _T_2503_0 <= _T_2503_1;
    _T_2503_1 <= io_inSprite_123;
    _T_2515_0 <= _T_2515_1;
    _T_2515_1 <= io_inSprite_124;
    _T_2527_0 <= _T_2527_1;
    _T_2527_1 <= io_inSprite_125;
    _T_2539_0 <= _T_2539_1;
    _T_2539_1 <= io_inSprite_126;
    _T_2551_0 <= _T_2551_1;
    _T_2551_1 <= io_inSprite_127;
  end
endmodule
module GraphicEngineVGA(
  input         clock,
  input         reset,
  input  [10:0] io_spriteXPosition_0,
  input  [10:0] io_spriteXPosition_1,
  input  [10:0] io_spriteXPosition_2,
  input  [10:0] io_spriteXPosition_3,
  input  [10:0] io_spriteXPosition_4,
  input  [10:0] io_spriteXPosition_5,
  input  [10:0] io_spriteXPosition_6,
  input  [10:0] io_spriteXPosition_7,
  input  [10:0] io_spriteXPosition_8,
  input  [10:0] io_spriteXPosition_9,
  input  [10:0] io_spriteXPosition_10,
  input  [10:0] io_spriteXPosition_11,
  input  [10:0] io_spriteXPosition_12,
  input  [10:0] io_spriteXPosition_13,
  input  [10:0] io_spriteXPosition_14,
  input  [10:0] io_spriteXPosition_15,
  input  [10:0] io_spriteXPosition_16,
  input  [10:0] io_spriteXPosition_17,
  input  [10:0] io_spriteXPosition_18,
  input  [10:0] io_spriteXPosition_19,
  input  [10:0] io_spriteXPosition_20,
  input  [10:0] io_spriteXPosition_21,
  input  [10:0] io_spriteXPosition_22,
  input  [10:0] io_spriteXPosition_23,
  input  [10:0] io_spriteXPosition_24,
  input  [10:0] io_spriteXPosition_25,
  input  [10:0] io_spriteXPosition_26,
  input  [10:0] io_spriteXPosition_27,
  input  [10:0] io_spriteXPosition_28,
  input  [10:0] io_spriteXPosition_29,
  input  [10:0] io_spriteXPosition_30,
  input  [10:0] io_spriteXPosition_31,
  input  [10:0] io_spriteXPosition_32,
  input  [10:0] io_spriteXPosition_33,
  input  [10:0] io_spriteXPosition_41,
  input  [10:0] io_spriteXPosition_42,
  input  [10:0] io_spriteXPosition_43,
  input  [10:0] io_spriteXPosition_44,
  input  [10:0] io_spriteXPosition_45,
  input  [10:0] io_spriteXPosition_46,
  input  [10:0] io_spriteXPosition_47,
  input  [10:0] io_spriteXPosition_48,
  input  [10:0] io_spriteXPosition_49,
  input  [10:0] io_spriteXPosition_50,
  input  [10:0] io_spriteXPosition_51,
  input  [10:0] io_spriteXPosition_122,
  input  [10:0] io_spriteXPosition_123,
  input  [10:0] io_spriteXPosition_124,
  input  [10:0] io_spriteXPosition_125,
  input  [10:0] io_spriteXPosition_126,
  input  [10:0] io_spriteXPosition_127,
  input  [9:0]  io_spriteYPosition_0,
  input  [9:0]  io_spriteYPosition_1,
  input  [9:0]  io_spriteYPosition_2,
  input  [9:0]  io_spriteYPosition_3,
  input  [9:0]  io_spriteYPosition_4,
  input  [9:0]  io_spriteYPosition_5,
  input  [9:0]  io_spriteYPosition_6,
  input  [9:0]  io_spriteYPosition_7,
  input  [9:0]  io_spriteYPosition_8,
  input  [9:0]  io_spriteYPosition_9,
  input  [9:0]  io_spriteYPosition_10,
  input  [9:0]  io_spriteYPosition_11,
  input  [9:0]  io_spriteYPosition_12,
  input  [9:0]  io_spriteYPosition_13,
  input  [9:0]  io_spriteYPosition_14,
  input  [9:0]  io_spriteYPosition_15,
  input  [9:0]  io_spriteYPosition_16,
  input  [9:0]  io_spriteYPosition_17,
  input  [9:0]  io_spriteYPosition_18,
  input  [9:0]  io_spriteYPosition_19,
  input  [9:0]  io_spriteYPosition_20,
  input  [9:0]  io_spriteYPosition_21,
  input  [9:0]  io_spriteYPosition_22,
  input  [9:0]  io_spriteYPosition_23,
  input  [9:0]  io_spriteYPosition_24,
  input  [9:0]  io_spriteYPosition_25,
  input  [9:0]  io_spriteYPosition_26,
  input  [9:0]  io_spriteYPosition_27,
  input  [9:0]  io_spriteYPosition_28,
  input  [9:0]  io_spriteYPosition_29,
  input  [9:0]  io_spriteYPosition_30,
  input  [9:0]  io_spriteYPosition_31,
  input  [9:0]  io_spriteYPosition_32,
  input  [9:0]  io_spriteYPosition_33,
  input  [9:0]  io_spriteYPosition_41,
  input  [9:0]  io_spriteYPosition_42,
  input  [9:0]  io_spriteYPosition_43,
  input  [9:0]  io_spriteYPosition_122,
  input  [9:0]  io_spriteYPosition_123,
  input  [9:0]  io_spriteYPosition_124,
  input  [9:0]  io_spriteYPosition_125,
  input  [9:0]  io_spriteYPosition_126,
  input  [9:0]  io_spriteYPosition_127,
  input         io_spriteVisible_0,
  input         io_spriteVisible_1,
  input         io_spriteVisible_2,
  input         io_spriteVisible_3,
  input         io_spriteVisible_4,
  input         io_spriteVisible_5,
  input         io_spriteVisible_6,
  input         io_spriteVisible_7,
  input         io_spriteVisible_8,
  input         io_spriteVisible_9,
  input         io_spriteVisible_10,
  input         io_spriteVisible_11,
  input         io_spriteVisible_12,
  input         io_spriteVisible_13,
  input         io_spriteVisible_14,
  input         io_spriteVisible_15,
  input         io_spriteVisible_16,
  input         io_spriteVisible_17,
  input         io_spriteVisible_18,
  input         io_spriteVisible_19,
  input         io_spriteVisible_20,
  input         io_spriteVisible_21,
  input         io_spriteVisible_22,
  input         io_spriteVisible_23,
  input         io_spriteVisible_24,
  input         io_spriteVisible_25,
  input         io_spriteVisible_26,
  input         io_spriteVisible_27,
  input         io_spriteVisible_28,
  input         io_spriteVisible_29,
  input         io_spriteVisible_30,
  input         io_spriteVisible_31,
  input         io_spriteVisible_32,
  input         io_spriteVisible_33,
  input         io_spriteVisible_41,
  input         io_spriteVisible_42,
  input         io_spriteVisible_43,
  input         io_spriteVisible_44,
  input         io_spriteVisible_45,
  input         io_spriteVisible_46,
  input         io_spriteVisible_47,
  input         io_spriteVisible_48,
  input         io_spriteVisible_49,
  input         io_spriteVisible_50,
  input         io_spriteVisible_51,
  input         io_spriteVisible_55,
  input         io_spriteVisible_56,
  input         io_spriteVisible_57,
  input         io_spriteVisible_61,
  input         io_spriteVisible_62,
  input         io_spriteVisible_63,
  input         io_spriteVisible_64,
  input         io_spriteVisible_65,
  input         io_spriteVisible_66,
  input         io_spriteVisible_70,
  input         io_spriteVisible_71,
  input         io_spriteVisible_72,
  input         io_spriteFlipVertical_122,
  input         io_spriteFlipVertical_123,
  input         io_spriteFlipVertical_124,
  input         io_spriteFlipVertical_125,
  input         io_spriteFlipVertical_126,
  input         io_spriteFlipVertical_127,
  input  [9:0]  io_viewBoxX_0,
  input  [4:0]  io_backBufferWriteData,
  input  [10:0] io_backBufferWriteAddress,
  input         io_backBufferWriteEnable,
  output        io_newFrame,
  input         io_frameUpdateDone,
  output        io_missingFrameError,
  output        io_backBufferWriteError,
  output        io_viewBoxOutOfRangeError,
  output [3:0]  io_vgaRed,
  output [3:0]  io_vgaBlue,
  output [3:0]  io_vgaGreen,
  output        io_Hsync,
  output        io_Vsync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
`endif // RANDOMIZE_REG_INIT
  wire  backTileMemories_0_0_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_0_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_0_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_1_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_1_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_1_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_2_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_2_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_2_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_3_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_3_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_3_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_4_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_4_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_4_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_5_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_5_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_5_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_6_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_6_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_6_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_7_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_7_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_7_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_8_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_8_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_8_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_9_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_9_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_9_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_10_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_10_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_10_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_11_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_11_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_11_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_12_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_12_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_12_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_13_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_13_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_13_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_14_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_14_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_14_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_15_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_15_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_15_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_16_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_16_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_16_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_17_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_17_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_17_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_18_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_18_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_18_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_19_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_19_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_19_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_20_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_20_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_20_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_21_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_21_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_21_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_22_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_22_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_22_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_23_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_23_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_23_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_24_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_24_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_24_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_25_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_25_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_25_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_26_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_26_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_26_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_27_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_27_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_27_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_28_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_28_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_28_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_29_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_29_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_29_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_30_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_30_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_30_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_0_31_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_0_31_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_0_31_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_0_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_0_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_0_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_1_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_1_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_1_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_2_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_2_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_2_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_3_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_3_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_3_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_4_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_4_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_4_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_5_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_5_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_5_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_6_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_6_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_6_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_7_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_7_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_7_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_8_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_8_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_8_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_9_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_9_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_9_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_10_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_10_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_10_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_11_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_11_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_11_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_12_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_12_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_12_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_13_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_13_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_13_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_14_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_14_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_14_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_15_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_15_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_15_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_16_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_16_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_16_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_17_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_17_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_17_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_18_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_18_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_18_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_19_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_19_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_19_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_20_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_20_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_20_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_21_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_21_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_21_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_22_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_22_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_22_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_23_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_23_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_23_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_24_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_24_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_24_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_25_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_25_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_25_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_26_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_26_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_26_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_27_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_27_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_27_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_28_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_28_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_28_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_29_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_29_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_29_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_30_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_30_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_30_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backTileMemories_1_31_clock; // @[GraphicEngineVGA.scala 205:34]
  wire [9:0] backTileMemories_1_31_io_address; // @[GraphicEngineVGA.scala 205:34]
  wire [6:0] backTileMemories_1_31_io_dataRead; // @[GraphicEngineVGA.scala 205:34]
  wire  backBufferMemories_0_clock; // @[GraphicEngineVGA.scala 230:34]
  wire [10:0] backBufferMemories_0_io_address; // @[GraphicEngineVGA.scala 230:34]
  wire [4:0] backBufferMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 230:34]
  wire  backBufferMemories_0_io_writeEnable; // @[GraphicEngineVGA.scala 230:34]
  wire [4:0] backBufferMemories_0_io_dataWrite; // @[GraphicEngineVGA.scala 230:34]
  wire  backBufferMemories_1_clock; // @[GraphicEngineVGA.scala 230:34]
  wire [10:0] backBufferMemories_1_io_address; // @[GraphicEngineVGA.scala 230:34]
  wire [4:0] backBufferMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 230:34]
  wire  backBufferMemories_1_io_writeEnable; // @[GraphicEngineVGA.scala 230:34]
  wire [4:0] backBufferMemories_1_io_dataWrite; // @[GraphicEngineVGA.scala 230:34]
  wire  backBufferShadowMemories_0_clock; // @[GraphicEngineVGA.scala 235:40]
  wire [10:0] backBufferShadowMemories_0_io_address; // @[GraphicEngineVGA.scala 235:40]
  wire [4:0] backBufferShadowMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 235:40]
  wire  backBufferShadowMemories_0_io_writeEnable; // @[GraphicEngineVGA.scala 235:40]
  wire [4:0] backBufferShadowMemories_0_io_dataWrite; // @[GraphicEngineVGA.scala 235:40]
  wire  backBufferShadowMemories_1_clock; // @[GraphicEngineVGA.scala 235:40]
  wire [10:0] backBufferShadowMemories_1_io_address; // @[GraphicEngineVGA.scala 235:40]
  wire [4:0] backBufferShadowMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 235:40]
  wire  backBufferShadowMemories_1_io_writeEnable; // @[GraphicEngineVGA.scala 235:40]
  wire [4:0] backBufferShadowMemories_1_io_dataWrite; // @[GraphicEngineVGA.scala 235:40]
  wire  backBufferRestoreMemories_0_clock; // @[GraphicEngineVGA.scala 241:41]
  wire [10:0] backBufferRestoreMemories_0_io_address; // @[GraphicEngineVGA.scala 241:41]
  wire [4:0] backBufferRestoreMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 241:41]
  wire  backBufferRestoreMemories_1_clock; // @[GraphicEngineVGA.scala 241:41]
  wire [10:0] backBufferRestoreMemories_1_io_address; // @[GraphicEngineVGA.scala 241:41]
  wire [4:0] backBufferRestoreMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 241:41]
  wire  spriteMemories_0_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_0_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_1_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_1_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_2_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_2_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_2_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_3_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_3_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_3_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_4_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_4_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_4_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_5_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_5_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_5_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_6_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_6_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_6_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_7_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_7_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_7_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_8_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_8_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_8_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_9_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_9_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_9_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_10_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_10_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_10_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_11_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_11_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_11_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_12_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_12_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_12_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_13_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_13_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_13_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_14_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_14_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_14_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_15_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_15_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_15_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_16_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_16_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_16_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_17_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_17_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_17_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_18_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_18_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_18_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_19_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_19_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_19_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_20_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_20_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_20_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_21_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_21_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_21_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_22_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_22_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_22_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_23_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_23_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_23_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_24_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_24_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_24_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_25_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_25_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_25_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_26_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_26_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_26_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_27_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_27_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_27_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_28_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_28_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_28_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_29_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_29_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_29_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_30_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_30_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_30_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_31_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_31_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_31_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_32_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_32_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_32_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_33_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_33_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_33_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_34_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_34_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_34_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_35_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_35_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_35_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_36_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_36_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_36_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_37_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_37_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_37_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_38_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_38_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_38_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_39_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_39_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_39_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_40_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_40_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_40_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_41_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_41_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_41_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_42_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_42_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_42_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_43_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_43_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_43_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_44_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_44_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_44_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_45_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_45_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_45_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_46_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_46_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_46_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_47_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_47_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_47_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_48_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_48_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_48_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_49_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_49_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_49_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_50_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_50_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_50_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_51_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_51_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_51_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_52_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_52_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_52_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_53_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_53_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_53_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_54_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_54_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_54_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_55_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_55_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_55_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_56_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_56_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_56_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_57_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_57_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_57_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_58_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_58_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_58_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_59_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_59_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_59_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_60_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_60_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_60_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_61_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_61_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_61_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_62_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_62_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_62_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_63_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_63_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_63_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_64_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_64_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_64_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_65_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_65_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_65_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_66_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_66_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_66_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_67_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_67_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_67_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_68_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_68_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_68_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_69_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_69_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_69_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_70_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_70_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_70_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_71_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_71_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_71_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_72_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_72_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_72_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_73_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_73_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_73_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_74_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_74_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_74_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_75_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_75_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_75_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_76_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_76_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_76_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_77_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_77_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_77_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_78_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_78_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_78_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_79_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_79_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_79_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_80_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_80_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_80_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_81_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_81_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_81_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_82_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_82_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_82_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_83_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_83_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_83_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_84_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_84_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_84_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_85_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_85_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_85_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_86_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_86_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_86_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_87_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_87_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_87_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_88_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_88_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_88_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_89_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_89_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_89_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_90_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_90_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_90_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_91_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_91_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_91_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_92_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_92_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_92_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_93_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_93_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_93_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_94_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_94_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_94_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_95_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_95_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_95_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_96_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_96_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_96_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_97_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_97_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_97_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_98_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_98_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_98_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_99_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_99_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_99_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_100_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_100_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_100_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_101_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_101_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_101_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_102_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_102_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_102_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_103_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_103_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_103_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_104_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_104_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_104_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_105_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_105_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_105_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_106_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_106_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_106_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_107_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_107_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_107_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_108_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_108_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_108_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_109_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_109_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_109_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_110_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_110_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_110_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_111_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_111_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_111_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_112_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_112_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_112_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_113_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_113_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_113_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_114_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_114_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_114_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_115_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_115_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_115_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_116_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_116_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_116_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_117_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_117_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_117_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_118_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_118_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_118_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_119_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_119_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_119_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_120_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_120_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_120_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_121_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_121_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_121_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_122_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_122_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_122_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_123_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_123_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_123_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_124_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_124_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_124_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_125_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_125_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_125_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_126_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_126_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_126_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  spriteMemories_127_clock; // @[GraphicEngineVGA.scala 320:30]
  wire [9:0] spriteMemories_127_io_address; // @[GraphicEngineVGA.scala 320:30]
  wire [6:0] spriteMemories_127_io_dataRead; // @[GraphicEngineVGA.scala 320:30]
  wire  rotation45deg_0_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_0_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_1_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_1_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_2_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_2_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_3_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_3_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_4_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_4_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_5_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_5_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_6_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_6_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_7_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_7_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_8_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_8_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_9_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_9_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_10_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_10_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_11_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_11_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_12_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_12_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_13_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_13_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_14_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_14_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_15_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_15_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_16_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_16_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_17_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_17_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_18_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_18_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_19_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_19_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_20_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_20_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_21_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_21_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_22_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_22_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_23_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_23_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_24_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_24_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_25_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_25_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_26_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_26_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_27_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_27_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_28_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_28_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_29_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_29_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_30_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_30_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_31_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_31_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_32_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_32_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_33_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_33_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_34_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_34_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_35_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_35_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_36_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_36_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_37_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_37_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_38_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_38_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_39_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_39_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_40_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_40_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_41_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_41_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_42_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_42_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_43_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_43_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_44_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_44_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_45_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_45_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_46_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_46_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_47_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_47_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_48_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_48_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_49_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_49_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_50_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_50_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_51_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_51_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_52_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_52_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_53_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_53_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_54_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_54_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_55_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_55_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_56_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_56_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_57_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_57_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_58_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_58_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_59_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_59_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_60_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_60_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_61_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_61_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_62_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_62_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_63_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_63_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_64_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_64_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_65_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_65_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_66_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_66_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_67_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_67_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_68_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_68_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_69_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_69_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_70_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_70_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_71_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_71_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_72_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_72_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_73_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_73_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_74_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_74_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_75_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_75_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_76_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_76_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_77_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_77_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_78_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_78_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_79_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_79_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_80_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_80_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_81_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_81_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_82_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_82_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_83_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_83_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_84_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_84_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_85_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_85_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_86_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_86_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_87_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_87_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_88_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_88_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_89_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_89_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_90_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_90_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_91_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_91_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_92_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_92_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_93_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_93_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_94_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_94_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_95_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_95_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_96_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_96_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_97_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_97_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_98_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_98_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_99_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_99_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_100_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_100_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_101_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_101_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_102_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_102_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_103_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_103_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_104_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_104_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_105_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_105_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_106_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_106_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_107_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_107_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_108_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_108_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_109_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_109_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_110_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_110_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_111_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_111_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_112_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_112_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_113_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_113_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_114_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_114_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_115_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_115_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_116_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_116_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_117_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_117_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_118_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_118_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_119_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_119_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_120_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_120_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_121_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_121_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_122_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_122_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_123_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_123_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_124_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_124_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_125_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_125_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_126_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_126_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  rotation45deg_127_clock; // @[GraphicEngineVGA.scala 325:30]
  wire [11:0] rotation45deg_127_io_address; // @[GraphicEngineVGA.scala 325:30]
  wire  spriteBlender_clock; // @[GraphicEngineVGA.scala 333:29]
  wire [5:0] spriteBlender_io_pixelColorBack; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_0; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_1; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_2; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_3; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_4; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_5; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_6; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_7; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_8; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_9; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_10; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_11; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_12; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_13; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_14; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_15; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_16; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_17; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_18; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_19; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_20; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_21; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_22; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_23; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_24; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_25; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_26; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_27; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_28; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_29; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_30; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_31; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_32; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_33; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_41; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_42; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_43; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_44; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_45; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_46; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_47; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_48; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_49; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_50; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_51; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_55; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_56; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_57; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_61; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_62; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_63; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_64; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_65; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_66; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_70; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_71; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_spriteVisibleReg_72; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_0; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_1; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_2; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_3; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_4; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_5; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_6; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_7; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_8; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_9; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_10; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_11; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_12; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_13; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_14; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_15; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_16; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_17; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_18; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_19; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_20; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_21; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_22; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_23; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_24; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_25; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_26; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_27; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_28; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_29; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_30; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_31; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_32; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_33; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_34; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_35; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_36; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_37; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_38; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_39; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_40; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_41; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_42; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_43; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_44; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_45; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_46; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_47; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_48; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_49; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_50; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_51; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_52; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_53; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_54; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_55; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_56; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_57; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_58; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_59; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_60; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_61; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_62; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_63; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_64; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_65; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_66; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_67; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_68; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_69; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_70; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_71; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_72; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_73; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_74; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_75; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_76; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_77; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_78; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_79; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_80; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_81; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_82; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_83; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_84; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_85; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_86; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_87; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_88; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_89; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_90; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_91; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_92; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_93; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_94; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_95; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_96; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_97; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_98; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_99; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_100; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_101; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_102; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_103; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_104; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_105; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_106; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_107; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_108; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_109; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_110; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_111; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_112; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_113; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_114; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_115; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_116; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_117; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_118; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_119; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_120; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_121; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_122; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_123; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_124; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_125; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_126; // @[GraphicEngineVGA.scala 333:29]
  wire  spriteBlender_io_inSprite_127; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_0; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_1; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_2; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_3; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_4; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_5; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_6; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_7; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_8; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_9; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_10; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_11; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_12; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_13; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_14; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_15; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_16; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_17; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_18; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_19; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_20; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_21; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_22; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_23; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_24; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_25; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_26; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_27; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_28; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_29; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_30; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_31; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_32; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_33; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_34; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_35; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_36; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_37; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_38; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_39; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_40; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_41; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_42; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_43; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_44; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_45; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_46; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_47; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_48; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_49; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_50; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_51; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_52; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_53; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_54; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_55; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_56; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_57; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_58; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_59; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_60; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_61; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_62; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_63; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_64; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_65; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_66; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_67; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_68; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_69; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_70; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_71; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_72; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_73; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_74; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_75; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_76; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_77; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_78; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_79; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_80; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_81; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_82; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_83; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_84; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_85; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_86; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_87; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_88; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_89; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_90; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_91; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_92; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_93; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_94; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_95; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_96; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_97; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_98; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_99; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_100; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_101; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_102; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_103; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_104; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_105; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_106; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_107; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_108; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_109; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_110; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_111; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_112; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_113; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_114; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_115; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_116; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_117; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_118; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_119; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_120; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_121; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_122; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_123; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_124; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_125; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_126; // @[GraphicEngineVGA.scala 333:29]
  wire [6:0] spriteBlender_io_datareader_127; // @[GraphicEngineVGA.scala 333:29]
  wire [3:0] spriteBlender_io_vgaRed; // @[GraphicEngineVGA.scala 333:29]
  wire [3:0] spriteBlender_io_vgaGreen; // @[GraphicEngineVGA.scala 333:29]
  wire [3:0] spriteBlender_io_vgaBlue; // @[GraphicEngineVGA.scala 333:29]
  reg [1:0] ScaleCounterReg; // @[GraphicEngineVGA.scala 73:32]
  reg [9:0] CounterXReg; // @[GraphicEngineVGA.scala 74:28]
  reg [9:0] CounterYReg; // @[GraphicEngineVGA.scala 75:28]
  wire  _T = ScaleCounterReg == 2'h3; // @[GraphicEngineVGA.scala 81:26]
  wire  _T_1 = CounterXReg == 10'h31f; // @[GraphicEngineVGA.scala 84:24]
  wire  _T_2 = CounterYReg == 10'h20c; // @[GraphicEngineVGA.scala 86:26]
  wire [9:0] _T_4 = CounterYReg + 10'h1; // @[GraphicEngineVGA.scala 90:38]
  wire [9:0] _T_6 = CounterXReg + 10'h1; // @[GraphicEngineVGA.scala 93:36]
  wire  _GEN_4 = _T_1 & _T_2; // @[GraphicEngineVGA.scala 84:129]
  wire [1:0] _T_8 = ScaleCounterReg + 2'h1; // @[GraphicEngineVGA.scala 96:42]
  wire  _GEN_8 = _T & _GEN_4; // @[GraphicEngineVGA.scala 81:52]
  reg [11:0] backMemoryRestoreCounter; // @[GraphicEngineVGA.scala 266:41]
  wire  restoreEnabled = backMemoryRestoreCounter < 12'h800; // @[GraphicEngineVGA.scala 269:33]
  wire  run = restoreEnabled ? 1'h0 : 1'h1; // @[GraphicEngineVGA.scala 269:70]
  wire  _T_9 = CounterXReg >= 10'h290; // @[GraphicEngineVGA.scala 100:28]
  wire  _T_10 = CounterXReg < 10'h2f0; // @[GraphicEngineVGA.scala 100:95]
  wire  Hsync = _T_9 & _T_10; // @[GraphicEngineVGA.scala 100:79]
  wire  _T_11 = CounterYReg >= 10'h1ea; // @[GraphicEngineVGA.scala 101:28]
  wire  _T_12 = CounterYReg < 10'h1ec; // @[GraphicEngineVGA.scala 101:95]
  wire  Vsync = _T_11 & _T_12; // @[GraphicEngineVGA.scala 101:79]
  reg  _T_14_0; // @[GameUtilities.scala 21:24]
  reg  _T_14_1; // @[GameUtilities.scala 21:24]
  reg  _T_14_2; // @[GameUtilities.scala 21:24]
  reg  _T_14_3; // @[GameUtilities.scala 21:24]
  reg  _T_16_0; // @[GameUtilities.scala 21:24]
  reg  _T_16_1; // @[GameUtilities.scala 21:24]
  reg  _T_16_2; // @[GameUtilities.scala 21:24]
  reg  _T_16_3; // @[GameUtilities.scala 21:24]
  wire  _T_17 = CounterXReg < 10'h280; // @[GraphicEngineVGA.scala 105:36]
  wire  _T_18 = CounterYReg < 10'h1e0; // @[GraphicEngineVGA.scala 105:76]
  reg [20:0] frameClockCount; // @[GraphicEngineVGA.scala 112:32]
  wire  _T_19 = frameClockCount == 21'h19a27f; // @[GraphicEngineVGA.scala 113:42]
  wire [20:0] _T_21 = frameClockCount + 21'h1; // @[GraphicEngineVGA.scala 113:92]
  wire  preDisplayArea = frameClockCount >= 21'h199a1b; // @[GraphicEngineVGA.scala 114:40]
  reg [10:0] spriteXPositionReg_0; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_1; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_2; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_3; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_4; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_5; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_6; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_7; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_8; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_9; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_10; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_11; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_12; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_13; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_14; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_15; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_16; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_17; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_18; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_19; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_20; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_21; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_22; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_23; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_24; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_25; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_26; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_27; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_28; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_29; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_30; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_31; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_32; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_33; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_34; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_35; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_36; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_37; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_38; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_39; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_40; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_41; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_42; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_43; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_44; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_45; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_46; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_47; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_48; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_49; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_50; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_51; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_52; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_53; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_54; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_55; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_56; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_57; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_58; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_59; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_60; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_61; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_62; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_63; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_64; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_65; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_66; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_67; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_68; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_69; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_70; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_71; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_72; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_73; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_74; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_75; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_76; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_77; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_78; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_79; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_80; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_81; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_82; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_83; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_84; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_85; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_86; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_87; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_88; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_89; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_90; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_91; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_92; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_93; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_94; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_95; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_96; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_97; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_98; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_99; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_100; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_101; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_102; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_103; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_104; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_105; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_106; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_107; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_108; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_109; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_110; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_111; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_112; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_113; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_114; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_115; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_116; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_117; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_118; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_119; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_120; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_121; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_122; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_123; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_124; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_125; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_126; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_127; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_0; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_1; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_2; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_3; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_4; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_5; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_6; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_7; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_8; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_9; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_10; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_11; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_12; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_13; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_14; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_15; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_16; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_17; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_18; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_19; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_20; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_21; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_22; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_23; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_24; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_25; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_26; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_27; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_28; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_29; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_30; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_31; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_32; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_33; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_34; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_35; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_36; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_37; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_38; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_39; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_40; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_41; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_42; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_43; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_44; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_45; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_46; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_47; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_48; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_49; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_50; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_51; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_52; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_53; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_54; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_55; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_56; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_57; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_58; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_59; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_60; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_61; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_62; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_63; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_70; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_71; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_72; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_73; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_74; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_75; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_76; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_77; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_78; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_79; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_80; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_81; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_82; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_83; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_84; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_85; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_86; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_87; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_88; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_89; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_90; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_91; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_92; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_93; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_94; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_95; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_96; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_97; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_98; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_99; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_100; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_101; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_102; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_103; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_104; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_105; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_106; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_107; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_108; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_109; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_110; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_111; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_112; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_113; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_114; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_115; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_116; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_117; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_118; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_119; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_120; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_121; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_122; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_123; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_124; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_125; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_126; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_127; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_0; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_1; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_2; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_3; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_4; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_5; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_6; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_7; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_8; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_9; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_10; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_11; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_12; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_13; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_14; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_15; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_16; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_17; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_18; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_19; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_20; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_21; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_22; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_23; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_24; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_25; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_26; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_27; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_28; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_29; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_30; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_31; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_32; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_33; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_41; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_42; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_43; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_44; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_45; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_46; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_47; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_48; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_49; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_50; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_51; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_55; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_56; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_57; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_61; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_62; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_63; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_64; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_65; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_66; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_70; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_71; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_72; // @[Reg.scala 27:20]
  wire  _GEN_269 = io_newFrame ? io_spriteVisible_0 : spriteVisibleReg_0; // @[Reg.scala 28:19]
  wire  _GEN_270 = io_newFrame ? io_spriteVisible_1 : spriteVisibleReg_1; // @[Reg.scala 28:19]
  wire  _GEN_271 = io_newFrame ? io_spriteVisible_2 : spriteVisibleReg_2; // @[Reg.scala 28:19]
  wire  _GEN_272 = io_newFrame ? io_spriteVisible_3 : spriteVisibleReg_3; // @[Reg.scala 28:19]
  wire  _GEN_273 = io_newFrame ? io_spriteVisible_4 : spriteVisibleReg_4; // @[Reg.scala 28:19]
  wire  _GEN_274 = io_newFrame ? io_spriteVisible_5 : spriteVisibleReg_5; // @[Reg.scala 28:19]
  wire  _GEN_275 = io_newFrame ? io_spriteVisible_6 : spriteVisibleReg_6; // @[Reg.scala 28:19]
  wire  _GEN_276 = io_newFrame ? io_spriteVisible_7 : spriteVisibleReg_7; // @[Reg.scala 28:19]
  wire  _GEN_277 = io_newFrame ? io_spriteVisible_8 : spriteVisibleReg_8; // @[Reg.scala 28:19]
  wire  _GEN_278 = io_newFrame ? io_spriteVisible_9 : spriteVisibleReg_9; // @[Reg.scala 28:19]
  wire  _GEN_279 = io_newFrame ? io_spriteVisible_10 : spriteVisibleReg_10; // @[Reg.scala 28:19]
  wire  _GEN_280 = io_newFrame ? io_spriteVisible_11 : spriteVisibleReg_11; // @[Reg.scala 28:19]
  wire  _GEN_281 = io_newFrame ? io_spriteVisible_12 : spriteVisibleReg_12; // @[Reg.scala 28:19]
  wire  _GEN_282 = io_newFrame ? io_spriteVisible_13 : spriteVisibleReg_13; // @[Reg.scala 28:19]
  wire  _GEN_283 = io_newFrame ? io_spriteVisible_14 : spriteVisibleReg_14; // @[Reg.scala 28:19]
  wire  _GEN_284 = io_newFrame ? io_spriteVisible_15 : spriteVisibleReg_15; // @[Reg.scala 28:19]
  wire  _GEN_285 = io_newFrame ? io_spriteVisible_16 : spriteVisibleReg_16; // @[Reg.scala 28:19]
  wire  _GEN_286 = io_newFrame ? io_spriteVisible_17 : spriteVisibleReg_17; // @[Reg.scala 28:19]
  wire  _GEN_287 = io_newFrame ? io_spriteVisible_18 : spriteVisibleReg_18; // @[Reg.scala 28:19]
  wire  _GEN_288 = io_newFrame ? io_spriteVisible_19 : spriteVisibleReg_19; // @[Reg.scala 28:19]
  wire  _GEN_289 = io_newFrame ? io_spriteVisible_20 : spriteVisibleReg_20; // @[Reg.scala 28:19]
  wire  _GEN_290 = io_newFrame ? io_spriteVisible_21 : spriteVisibleReg_21; // @[Reg.scala 28:19]
  wire  _GEN_291 = io_newFrame ? io_spriteVisible_22 : spriteVisibleReg_22; // @[Reg.scala 28:19]
  wire  _GEN_292 = io_newFrame ? io_spriteVisible_23 : spriteVisibleReg_23; // @[Reg.scala 28:19]
  wire  _GEN_293 = io_newFrame ? io_spriteVisible_24 : spriteVisibleReg_24; // @[Reg.scala 28:19]
  wire  _GEN_294 = io_newFrame ? io_spriteVisible_25 : spriteVisibleReg_25; // @[Reg.scala 28:19]
  wire  _GEN_295 = io_newFrame ? io_spriteVisible_26 : spriteVisibleReg_26; // @[Reg.scala 28:19]
  wire  _GEN_296 = io_newFrame ? io_spriteVisible_27 : spriteVisibleReg_27; // @[Reg.scala 28:19]
  wire  _GEN_297 = io_newFrame ? io_spriteVisible_28 : spriteVisibleReg_28; // @[Reg.scala 28:19]
  wire  _GEN_298 = io_newFrame ? io_spriteVisible_29 : spriteVisibleReg_29; // @[Reg.scala 28:19]
  wire  _GEN_299 = io_newFrame ? io_spriteVisible_30 : spriteVisibleReg_30; // @[Reg.scala 28:19]
  wire  _GEN_300 = io_newFrame ? io_spriteVisible_31 : spriteVisibleReg_31; // @[Reg.scala 28:19]
  wire  _GEN_301 = io_newFrame ? io_spriteVisible_32 : spriteVisibleReg_32; // @[Reg.scala 28:19]
  wire  _GEN_302 = io_newFrame ? io_spriteVisible_33 : spriteVisibleReg_33; // @[Reg.scala 28:19]
  wire  _GEN_310 = io_newFrame ? io_spriteVisible_41 : spriteVisibleReg_41; // @[Reg.scala 28:19]
  wire  _GEN_311 = io_newFrame ? io_spriteVisible_42 : spriteVisibleReg_42; // @[Reg.scala 28:19]
  wire  _GEN_312 = io_newFrame ? io_spriteVisible_43 : spriteVisibleReg_43; // @[Reg.scala 28:19]
  wire  _GEN_313 = io_newFrame ? io_spriteVisible_44 : spriteVisibleReg_44; // @[Reg.scala 28:19]
  wire  _GEN_314 = io_newFrame ? io_spriteVisible_45 : spriteVisibleReg_45; // @[Reg.scala 28:19]
  wire  _GEN_315 = io_newFrame ? io_spriteVisible_46 : spriteVisibleReg_46; // @[Reg.scala 28:19]
  wire  _GEN_316 = io_newFrame ? io_spriteVisible_47 : spriteVisibleReg_47; // @[Reg.scala 28:19]
  wire  _GEN_317 = io_newFrame ? io_spriteVisible_48 : spriteVisibleReg_48; // @[Reg.scala 28:19]
  wire  _GEN_318 = io_newFrame ? io_spriteVisible_49 : spriteVisibleReg_49; // @[Reg.scala 28:19]
  wire  _GEN_319 = io_newFrame ? io_spriteVisible_50 : spriteVisibleReg_50; // @[Reg.scala 28:19]
  wire  _GEN_320 = io_newFrame ? io_spriteVisible_51 : spriteVisibleReg_51; // @[Reg.scala 28:19]
  wire  _GEN_324 = io_newFrame ? io_spriteVisible_55 : spriteVisibleReg_55; // @[Reg.scala 28:19]
  wire  _GEN_325 = io_newFrame ? io_spriteVisible_56 : spriteVisibleReg_56; // @[Reg.scala 28:19]
  wire  _GEN_326 = io_newFrame ? io_spriteVisible_57 : spriteVisibleReg_57; // @[Reg.scala 28:19]
  wire  _GEN_330 = io_newFrame ? io_spriteVisible_61 : spriteVisibleReg_61; // @[Reg.scala 28:19]
  wire  _GEN_331 = io_newFrame ? io_spriteVisible_62 : spriteVisibleReg_62; // @[Reg.scala 28:19]
  wire  _GEN_332 = io_newFrame ? io_spriteVisible_63 : spriteVisibleReg_63; // @[Reg.scala 28:19]
  wire  _GEN_333 = io_newFrame ? io_spriteVisible_64 : spriteVisibleReg_64; // @[Reg.scala 28:19]
  wire  _GEN_334 = io_newFrame ? io_spriteVisible_65 : spriteVisibleReg_65; // @[Reg.scala 28:19]
  wire  _GEN_335 = io_newFrame ? io_spriteVisible_66 : spriteVisibleReg_66; // @[Reg.scala 28:19]
  wire  _GEN_339 = io_newFrame ? io_spriteVisible_70 : spriteVisibleReg_70; // @[Reg.scala 28:19]
  wire  _GEN_340 = io_newFrame ? io_spriteVisible_71 : spriteVisibleReg_71; // @[Reg.scala 28:19]
  wire  _GEN_341 = io_newFrame ? io_spriteVisible_72 : spriteVisibleReg_72; // @[Reg.scala 28:19]
  reg  spriteFlipVerticalReg_122; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_123; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_124; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_125; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_126; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_127; // @[Reg.scala 27:20]
  reg [9:0] viewBoxXReg_0; // @[Reg.scala 27:20]
  reg  missingFrameErrorReg; // @[GraphicEngineVGA.scala 146:37]
  reg  backBufferWriteErrorReg; // @[GraphicEngineVGA.scala 147:40]
  reg  viewBoxOutOfRangeErrorReg; // @[GraphicEngineVGA.scala 148:42]
  wire  _T_32 = viewBoxXReg_0 >= 10'h280; // @[GraphicEngineVGA.scala 166:45]
  wire [9:0] viewBoxXClipped_0 = _T_32 ? 10'h280 : viewBoxXReg_0; // @[GraphicEngineVGA.scala 166:29]
  wire [10:0] pixelXBack_0 = CounterXReg + viewBoxXClipped_0; // @[GraphicEngineVGA.scala 168:29]
  wire [10:0] pixelYBack_0 = {{1'd0}, CounterYReg}; // @[GraphicEngineVGA.scala 169:29]
  wire [10:0] pixelXBack_1 = {{1'd0}, CounterXReg}; // @[GraphicEngineVGA.scala 168:29]
  wire  _T_44 = viewBoxXReg_0 > 10'h280; // @[GraphicEngineVGA.scala 172:23]
  wire  _GEN_1169 = _T_44 | viewBoxOutOfRangeErrorReg; // @[GraphicEngineVGA.scala 172:58]
  reg  newFrameStikyReg; // @[GraphicEngineVGA.scala 178:33]
  wire  _GEN_1170 = io_newFrame | newFrameStikyReg; // @[GraphicEngineVGA.scala 179:21]
  reg  _T_47; // @[GraphicEngineVGA.scala 182:15]
  wire  _T_48 = newFrameStikyReg & io_newFrame; // @[GraphicEngineVGA.scala 185:25]
  wire  _GEN_1172 = _T_48 | missingFrameErrorReg; // @[GraphicEngineVGA.scala 185:41]
  wire [5:0] _GEN_1246 = {{1'd0}, pixelYBack_0[4:0]}; // @[GraphicEngineVGA.scala 220:82]
  wire [10:0] _T_51 = 6'h20 * _GEN_1246; // @[GraphicEngineVGA.scala 220:82]
  wire [10:0] _GEN_1247 = {{6'd0}, pixelXBack_0[4:0]}; // @[GraphicEngineVGA.scala 220:69]
  wire [11:0] _T_52 = _GEN_1247 + _T_51; // @[GraphicEngineVGA.scala 220:69]
  reg [6:0] backTileMemoryDataRead_0_0; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_1; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_2; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_3; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_4; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_5; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_6; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_7; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_8; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_9; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_10; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_11; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_12; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_13; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_14; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_15; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_16; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_17; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_18; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_19; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_20; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_21; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_22; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_23; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_24; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_25; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_26; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_27; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_28; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_29; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_30; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_0_31; // @[GraphicEngineVGA.scala 222:44]
  wire [10:0] _GEN_1311 = {{6'd0}, pixelXBack_1[4:0]}; // @[GraphicEngineVGA.scala 220:69]
  wire [11:0] _T_212 = _GEN_1311 + _T_51; // @[GraphicEngineVGA.scala 220:69]
  reg [6:0] backTileMemoryDataRead_1_0; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_1; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_2; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_3; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_4; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_5; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_6; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_7; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_8; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_9; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_10; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_11; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_12; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_13; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_14; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_15; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_16; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_17; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_18; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_19; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_20; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_21; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_22; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_23; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_24; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_25; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_26; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_27; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_28; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_29; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_30; // @[GraphicEngineVGA.scala 222:44]
  reg [6:0] backTileMemoryDataRead_1_31; // @[GraphicEngineVGA.scala 222:44]
  reg [11:0] backMemoryCopyCounter; // @[GraphicEngineVGA.scala 247:38]
  wire  _T_369 = backMemoryCopyCounter < 12'h800; // @[GraphicEngineVGA.scala 251:32]
  wire [11:0] _T_371 = backMemoryCopyCounter + 12'h1; // @[GraphicEngineVGA.scala 252:54]
  wire  copyEnabled = preDisplayArea & _T_369; // @[GraphicEngineVGA.scala 250:24]
  reg  copyEnabledReg; // @[GraphicEngineVGA.scala 264:31]
  wire [11:0] _T_374 = backMemoryRestoreCounter + 12'h1; // @[GraphicEngineVGA.scala 270:58]
  reg [10:0] _T_377; // @[GraphicEngineVGA.scala 287:72]
  reg [10:0] _T_379; // @[GraphicEngineVGA.scala 287:161]
  wire [10:0] _T_380 = copyEnabled ? backMemoryCopyCounter[10:0] : _T_379; // @[GraphicEngineVGA.scala 287:110]
  reg  _T_382; // @[GraphicEngineVGA.scala 289:76]
  reg  _T_383; // @[GraphicEngineVGA.scala 289:127]
  wire  _T_384 = copyEnabled ? 1'h0 : _T_383; // @[GraphicEngineVGA.scala 289:97]
  reg [4:0] _T_386; // @[GraphicEngineVGA.scala 290:116]
  reg [10:0] _T_389; // @[GraphicEngineVGA.scala 292:66]
  wire [11:0] _T_392 = 6'h28 * pixelYBack_0[10:5]; // @[GraphicEngineVGA.scala 292:139]
  wire [11:0] _GEN_1374 = {{6'd0}, pixelXBack_0[10:5]}; // @[GraphicEngineVGA.scala 292:126]
  wire [12:0] _T_393 = _GEN_1374 + _T_392; // @[GraphicEngineVGA.scala 292:126]
  wire [12:0] _T_394 = copyEnabledReg ? {{2'd0}, _T_389} : _T_393; // @[GraphicEngineVGA.scala 292:42]
  reg [10:0] _T_397; // @[GraphicEngineVGA.scala 287:72]
  reg [10:0] _T_399; // @[GraphicEngineVGA.scala 287:161]
  wire [10:0] _T_400 = copyEnabled ? backMemoryCopyCounter[10:0] : _T_399; // @[GraphicEngineVGA.scala 287:110]
  reg  _T_402; // @[GraphicEngineVGA.scala 289:76]
  reg  _T_403; // @[GraphicEngineVGA.scala 289:127]
  wire  _T_404 = copyEnabled ? 1'h0 : _T_403; // @[GraphicEngineVGA.scala 289:97]
  reg [4:0] _T_406; // @[GraphicEngineVGA.scala 290:116]
  reg [10:0] _T_409; // @[GraphicEngineVGA.scala 292:66]
  wire [11:0] _GEN_1375 = {{6'd0}, pixelXBack_1[10:5]}; // @[GraphicEngineVGA.scala 292:126]
  wire [12:0] _T_413 = _GEN_1375 + _T_392; // @[GraphicEngineVGA.scala 292:126]
  wire [12:0] _T_414 = copyEnabledReg ? {{2'd0}, _T_409} : _T_413; // @[GraphicEngineVGA.scala 292:42]
  wire  _T_415 = copyEnabled | copyEnabledReg; // @[GraphicEngineVGA.scala 300:20]
  wire  _GEN_1180 = io_backBufferWriteEnable | backBufferWriteErrorReg; // @[GraphicEngineVGA.scala 301:36]
  reg [4:0] _T_416; // @[GraphicEngineVGA.scala 311:64]
  wire [6:0] _GEN_1183 = 5'h1 == _T_416 ? backTileMemoryDataRead_0_1 : backTileMemoryDataRead_0_0; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1184 = 5'h2 == _T_416 ? backTileMemoryDataRead_0_2 : _GEN_1183; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1185 = 5'h3 == _T_416 ? backTileMemoryDataRead_0_3 : _GEN_1184; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1186 = 5'h4 == _T_416 ? backTileMemoryDataRead_0_4 : _GEN_1185; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1187 = 5'h5 == _T_416 ? backTileMemoryDataRead_0_5 : _GEN_1186; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1188 = 5'h6 == _T_416 ? backTileMemoryDataRead_0_6 : _GEN_1187; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1189 = 5'h7 == _T_416 ? backTileMemoryDataRead_0_7 : _GEN_1188; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1190 = 5'h8 == _T_416 ? backTileMemoryDataRead_0_8 : _GEN_1189; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1191 = 5'h9 == _T_416 ? backTileMemoryDataRead_0_9 : _GEN_1190; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1192 = 5'ha == _T_416 ? backTileMemoryDataRead_0_10 : _GEN_1191; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1193 = 5'hb == _T_416 ? backTileMemoryDataRead_0_11 : _GEN_1192; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1194 = 5'hc == _T_416 ? backTileMemoryDataRead_0_12 : _GEN_1193; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1195 = 5'hd == _T_416 ? backTileMemoryDataRead_0_13 : _GEN_1194; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1196 = 5'he == _T_416 ? backTileMemoryDataRead_0_14 : _GEN_1195; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1197 = 5'hf == _T_416 ? backTileMemoryDataRead_0_15 : _GEN_1196; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1198 = 5'h10 == _T_416 ? backTileMemoryDataRead_0_16 : _GEN_1197; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1199 = 5'h11 == _T_416 ? backTileMemoryDataRead_0_17 : _GEN_1198; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1200 = 5'h12 == _T_416 ? backTileMemoryDataRead_0_18 : _GEN_1199; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1201 = 5'h13 == _T_416 ? backTileMemoryDataRead_0_19 : _GEN_1200; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1202 = 5'h14 == _T_416 ? backTileMemoryDataRead_0_20 : _GEN_1201; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1203 = 5'h15 == _T_416 ? backTileMemoryDataRead_0_21 : _GEN_1202; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1204 = 5'h16 == _T_416 ? backTileMemoryDataRead_0_22 : _GEN_1203; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1205 = 5'h17 == _T_416 ? backTileMemoryDataRead_0_23 : _GEN_1204; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1206 = 5'h18 == _T_416 ? backTileMemoryDataRead_0_24 : _GEN_1205; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1207 = 5'h19 == _T_416 ? backTileMemoryDataRead_0_25 : _GEN_1206; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1208 = 5'h1a == _T_416 ? backTileMemoryDataRead_0_26 : _GEN_1207; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1209 = 5'h1b == _T_416 ? backTileMemoryDataRead_0_27 : _GEN_1208; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1210 = 5'h1c == _T_416 ? backTileMemoryDataRead_0_28 : _GEN_1209; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1211 = 5'h1d == _T_416 ? backTileMemoryDataRead_0_29 : _GEN_1210; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1212 = 5'h1e == _T_416 ? backTileMemoryDataRead_0_30 : _GEN_1211; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] fullBackgroundColor_0 = 5'h1f == _T_416 ? backTileMemoryDataRead_0_31 : _GEN_1212; // @[GraphicEngineVGA.scala 311:28]
  reg [4:0] _T_419; // @[GraphicEngineVGA.scala 311:64]
  wire [6:0] _GEN_1215 = 5'h1 == _T_419 ? backTileMemoryDataRead_1_1 : backTileMemoryDataRead_1_0; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1216 = 5'h2 == _T_419 ? backTileMemoryDataRead_1_2 : _GEN_1215; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1217 = 5'h3 == _T_419 ? backTileMemoryDataRead_1_3 : _GEN_1216; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1218 = 5'h4 == _T_419 ? backTileMemoryDataRead_1_4 : _GEN_1217; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1219 = 5'h5 == _T_419 ? backTileMemoryDataRead_1_5 : _GEN_1218; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1220 = 5'h6 == _T_419 ? backTileMemoryDataRead_1_6 : _GEN_1219; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1221 = 5'h7 == _T_419 ? backTileMemoryDataRead_1_7 : _GEN_1220; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1222 = 5'h8 == _T_419 ? backTileMemoryDataRead_1_8 : _GEN_1221; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1223 = 5'h9 == _T_419 ? backTileMemoryDataRead_1_9 : _GEN_1222; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1224 = 5'ha == _T_419 ? backTileMemoryDataRead_1_10 : _GEN_1223; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1225 = 5'hb == _T_419 ? backTileMemoryDataRead_1_11 : _GEN_1224; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1226 = 5'hc == _T_419 ? backTileMemoryDataRead_1_12 : _GEN_1225; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1227 = 5'hd == _T_419 ? backTileMemoryDataRead_1_13 : _GEN_1226; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1228 = 5'he == _T_419 ? backTileMemoryDataRead_1_14 : _GEN_1227; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1229 = 5'hf == _T_419 ? backTileMemoryDataRead_1_15 : _GEN_1228; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1230 = 5'h10 == _T_419 ? backTileMemoryDataRead_1_16 : _GEN_1229; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1231 = 5'h11 == _T_419 ? backTileMemoryDataRead_1_17 : _GEN_1230; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1232 = 5'h12 == _T_419 ? backTileMemoryDataRead_1_18 : _GEN_1231; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1233 = 5'h13 == _T_419 ? backTileMemoryDataRead_1_19 : _GEN_1232; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1234 = 5'h14 == _T_419 ? backTileMemoryDataRead_1_20 : _GEN_1233; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1235 = 5'h15 == _T_419 ? backTileMemoryDataRead_1_21 : _GEN_1234; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1236 = 5'h16 == _T_419 ? backTileMemoryDataRead_1_22 : _GEN_1235; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1237 = 5'h17 == _T_419 ? backTileMemoryDataRead_1_23 : _GEN_1236; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1238 = 5'h18 == _T_419 ? backTileMemoryDataRead_1_24 : _GEN_1237; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1239 = 5'h19 == _T_419 ? backTileMemoryDataRead_1_25 : _GEN_1238; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1240 = 5'h1a == _T_419 ? backTileMemoryDataRead_1_26 : _GEN_1239; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1241 = 5'h1b == _T_419 ? backTileMemoryDataRead_1_27 : _GEN_1240; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1242 = 5'h1c == _T_419 ? backTileMemoryDataRead_1_28 : _GEN_1241; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1243 = 5'h1d == _T_419 ? backTileMemoryDataRead_1_29 : _GEN_1242; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] _GEN_1244 = 5'h1e == _T_419 ? backTileMemoryDataRead_1_30 : _GEN_1243; // @[GraphicEngineVGA.scala 311:28]
  wire [6:0] fullBackgroundColor_1 = 5'h1f == _T_419 ? backTileMemoryDataRead_1_31 : _GEN_1244; // @[GraphicEngineVGA.scala 311:28]
  reg [5:0] pixelColorBack; // @[GraphicEngineVGA.scala 314:31]
  wire [10:0] _T_438 = {1'h0,CounterXReg}; // @[GraphicEngineVGA.scala 355:52]
  reg [11:0] inSpriteX_0; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _T_442 = {1'h0,CounterYReg}; // @[GraphicEngineVGA.scala 356:52]
  wire [10:0] _GEN_1376 = {{1{spriteYPositionReg_0[9]}},spriteYPositionReg_0}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_444; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_0 = _T_444[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [7:0] _T_464 = 8'sh20 - 8'sh1; // @[GraphicEngineVGA.scala 370:52]
  wire [11:0] _GEN_1378 = {{4{_T_464[7]}},_T_464}; // @[GraphicEngineVGA.scala 370:60]
  wire [11:0] _T_468 = {{1{inSpriteY_0[10]}},inSpriteY_0}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_486 = inSpriteX_0; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_494 = {{2'd0}, _T_486}; // @[Mux.scala 80:57]
  wire [11:0] _T_498 = {{1{inSpriteY_0[10]}},inSpriteY_0}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_506 = {{2'd0}, _T_498}; // @[Mux.scala 80:57]
  wire  _T_507 = $signed(inSpriteX_0) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_508 = $signed(inSpriteX_0) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_509 = _T_507 & _T_508; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_510 = $signed(_T_468) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_511 = $signed(_T_468) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_512 = _T_510 & _T_511; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_535 = _T_506 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1382 = {{7'd0}, _T_494}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_537 = _T_535 + _GEN_1382; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_1; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1385 = {{1{spriteYPositionReg_1[9]}},spriteYPositionReg_1}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_563; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_1 = _T_563[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_587 = {{1{inSpriteY_1[10]}},inSpriteY_1}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_605 = inSpriteX_1; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_613 = {{2'd0}, _T_605}; // @[Mux.scala 80:57]
  wire [11:0] _T_617 = {{1{inSpriteY_1[10]}},inSpriteY_1}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_625 = {{2'd0}, _T_617}; // @[Mux.scala 80:57]
  wire  _T_626 = $signed(inSpriteX_1) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_627 = $signed(inSpriteX_1) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_628 = _T_626 & _T_627; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_629 = $signed(_T_587) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_630 = $signed(_T_587) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_631 = _T_629 & _T_630; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_654 = _T_625 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1391 = {{7'd0}, _T_613}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_656 = _T_654 + _GEN_1391; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_2; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1394 = {{1{spriteYPositionReg_2[9]}},spriteYPositionReg_2}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_682; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_2 = _T_682[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_706 = {{1{inSpriteY_2[10]}},inSpriteY_2}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_724 = inSpriteX_2; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_732 = {{2'd0}, _T_724}; // @[Mux.scala 80:57]
  wire [11:0] _T_736 = {{1{inSpriteY_2[10]}},inSpriteY_2}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_744 = {{2'd0}, _T_736}; // @[Mux.scala 80:57]
  wire  _T_745 = $signed(inSpriteX_2) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_746 = $signed(inSpriteX_2) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_747 = _T_745 & _T_746; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_748 = $signed(_T_706) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_749 = $signed(_T_706) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_750 = _T_748 & _T_749; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_773 = _T_744 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1400 = {{7'd0}, _T_732}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_775 = _T_773 + _GEN_1400; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_3; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1403 = {{1{spriteYPositionReg_3[9]}},spriteYPositionReg_3}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_801; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_3 = _T_801[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_825 = {{1{inSpriteY_3[10]}},inSpriteY_3}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_843 = inSpriteX_3; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_851 = {{2'd0}, _T_843}; // @[Mux.scala 80:57]
  wire [11:0] _T_855 = {{1{inSpriteY_3[10]}},inSpriteY_3}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_863 = {{2'd0}, _T_855}; // @[Mux.scala 80:57]
  wire  _T_864 = $signed(inSpriteX_3) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_865 = $signed(inSpriteX_3) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_866 = _T_864 & _T_865; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_867 = $signed(_T_825) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_868 = $signed(_T_825) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_869 = _T_867 & _T_868; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_892 = _T_863 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1409 = {{7'd0}, _T_851}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_894 = _T_892 + _GEN_1409; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_4; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1412 = {{1{spriteYPositionReg_4[9]}},spriteYPositionReg_4}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_920; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_4 = _T_920[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_944 = {{1{inSpriteY_4[10]}},inSpriteY_4}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_962 = inSpriteX_4; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_970 = {{2'd0}, _T_962}; // @[Mux.scala 80:57]
  wire [11:0] _T_974 = {{1{inSpriteY_4[10]}},inSpriteY_4}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_982 = {{2'd0}, _T_974}; // @[Mux.scala 80:57]
  wire  _T_983 = $signed(inSpriteX_4) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_984 = $signed(inSpriteX_4) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_985 = _T_983 & _T_984; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_986 = $signed(_T_944) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_987 = $signed(_T_944) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_988 = _T_986 & _T_987; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1011 = _T_982 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1418 = {{7'd0}, _T_970}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1013 = _T_1011 + _GEN_1418; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_5; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1421 = {{1{spriteYPositionReg_5[9]}},spriteYPositionReg_5}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1039; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_5 = _T_1039[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1063 = {{1{inSpriteY_5[10]}},inSpriteY_5}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1081 = inSpriteX_5; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1089 = {{2'd0}, _T_1081}; // @[Mux.scala 80:57]
  wire [11:0] _T_1093 = {{1{inSpriteY_5[10]}},inSpriteY_5}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1101 = {{2'd0}, _T_1093}; // @[Mux.scala 80:57]
  wire  _T_1102 = $signed(inSpriteX_5) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1103 = $signed(inSpriteX_5) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1104 = _T_1102 & _T_1103; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1105 = $signed(_T_1063) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1106 = $signed(_T_1063) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1107 = _T_1105 & _T_1106; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1130 = _T_1101 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1427 = {{7'd0}, _T_1089}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1132 = _T_1130 + _GEN_1427; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_6; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1430 = {{1{spriteYPositionReg_6[9]}},spriteYPositionReg_6}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1158; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_6 = _T_1158[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1182 = {{1{inSpriteY_6[10]}},inSpriteY_6}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1200 = inSpriteX_6; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1208 = {{2'd0}, _T_1200}; // @[Mux.scala 80:57]
  wire [11:0] _T_1212 = {{1{inSpriteY_6[10]}},inSpriteY_6}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1220 = {{2'd0}, _T_1212}; // @[Mux.scala 80:57]
  wire  _T_1221 = $signed(inSpriteX_6) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1222 = $signed(inSpriteX_6) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1223 = _T_1221 & _T_1222; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1224 = $signed(_T_1182) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1225 = $signed(_T_1182) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1226 = _T_1224 & _T_1225; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1249 = _T_1220 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1436 = {{7'd0}, _T_1208}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1251 = _T_1249 + _GEN_1436; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_7; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1439 = {{1{spriteYPositionReg_7[9]}},spriteYPositionReg_7}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1277; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_7 = _T_1277[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1301 = {{1{inSpriteY_7[10]}},inSpriteY_7}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1319 = inSpriteX_7; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1327 = {{2'd0}, _T_1319}; // @[Mux.scala 80:57]
  wire [11:0] _T_1331 = {{1{inSpriteY_7[10]}},inSpriteY_7}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1339 = {{2'd0}, _T_1331}; // @[Mux.scala 80:57]
  wire  _T_1340 = $signed(inSpriteX_7) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1341 = $signed(inSpriteX_7) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1342 = _T_1340 & _T_1341; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1343 = $signed(_T_1301) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1344 = $signed(_T_1301) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1345 = _T_1343 & _T_1344; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1368 = _T_1339 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1445 = {{7'd0}, _T_1327}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1370 = _T_1368 + _GEN_1445; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_8; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1448 = {{1{spriteYPositionReg_8[9]}},spriteYPositionReg_8}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1396; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_8 = _T_1396[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1420 = {{1{inSpriteY_8[10]}},inSpriteY_8}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1438 = inSpriteX_8; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1446 = {{2'd0}, _T_1438}; // @[Mux.scala 80:57]
  wire [11:0] _T_1450 = {{1{inSpriteY_8[10]}},inSpriteY_8}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1458 = {{2'd0}, _T_1450}; // @[Mux.scala 80:57]
  wire  _T_1459 = $signed(inSpriteX_8) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1460 = $signed(inSpriteX_8) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1461 = _T_1459 & _T_1460; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1462 = $signed(_T_1420) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1463 = $signed(_T_1420) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1464 = _T_1462 & _T_1463; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1487 = _T_1458 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1454 = {{7'd0}, _T_1446}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1489 = _T_1487 + _GEN_1454; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_9; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1457 = {{1{spriteYPositionReg_9[9]}},spriteYPositionReg_9}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1515; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_9 = _T_1515[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1539 = {{1{inSpriteY_9[10]}},inSpriteY_9}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1557 = inSpriteX_9; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1565 = {{2'd0}, _T_1557}; // @[Mux.scala 80:57]
  wire [11:0] _T_1569 = {{1{inSpriteY_9[10]}},inSpriteY_9}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1577 = {{2'd0}, _T_1569}; // @[Mux.scala 80:57]
  wire  _T_1578 = $signed(inSpriteX_9) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1579 = $signed(inSpriteX_9) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1580 = _T_1578 & _T_1579; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1581 = $signed(_T_1539) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1582 = $signed(_T_1539) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1583 = _T_1581 & _T_1582; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1606 = _T_1577 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1463 = {{7'd0}, _T_1565}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1608 = _T_1606 + _GEN_1463; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_10; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1466 = {{1{spriteYPositionReg_10[9]}},spriteYPositionReg_10}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1634; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_10 = _T_1634[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1658 = {{1{inSpriteY_10[10]}},inSpriteY_10}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1676 = inSpriteX_10; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1684 = {{2'd0}, _T_1676}; // @[Mux.scala 80:57]
  wire [11:0] _T_1688 = {{1{inSpriteY_10[10]}},inSpriteY_10}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1696 = {{2'd0}, _T_1688}; // @[Mux.scala 80:57]
  wire  _T_1697 = $signed(inSpriteX_10) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1698 = $signed(inSpriteX_10) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1699 = _T_1697 & _T_1698; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1700 = $signed(_T_1658) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1701 = $signed(_T_1658) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1702 = _T_1700 & _T_1701; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1725 = _T_1696 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1472 = {{7'd0}, _T_1684}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1727 = _T_1725 + _GEN_1472; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_11; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1475 = {{1{spriteYPositionReg_11[9]}},spriteYPositionReg_11}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1753; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_11 = _T_1753[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1777 = {{1{inSpriteY_11[10]}},inSpriteY_11}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1795 = inSpriteX_11; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1803 = {{2'd0}, _T_1795}; // @[Mux.scala 80:57]
  wire [11:0] _T_1807 = {{1{inSpriteY_11[10]}},inSpriteY_11}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1815 = {{2'd0}, _T_1807}; // @[Mux.scala 80:57]
  wire  _T_1816 = $signed(inSpriteX_11) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1817 = $signed(inSpriteX_11) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1818 = _T_1816 & _T_1817; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1819 = $signed(_T_1777) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1820 = $signed(_T_1777) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1821 = _T_1819 & _T_1820; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1844 = _T_1815 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1481 = {{7'd0}, _T_1803}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1846 = _T_1844 + _GEN_1481; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_12; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1484 = {{1{spriteYPositionReg_12[9]}},spriteYPositionReg_12}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1872; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_12 = _T_1872[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_1896 = {{1{inSpriteY_12[10]}},inSpriteY_12}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_1914 = inSpriteX_12; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_1922 = {{2'd0}, _T_1914}; // @[Mux.scala 80:57]
  wire [11:0] _T_1926 = {{1{inSpriteY_12[10]}},inSpriteY_12}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_1934 = {{2'd0}, _T_1926}; // @[Mux.scala 80:57]
  wire  _T_1935 = $signed(inSpriteX_12) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_1936 = $signed(inSpriteX_12) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_1937 = _T_1935 & _T_1936; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_1938 = $signed(_T_1896) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_1939 = $signed(_T_1896) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_1940 = _T_1938 & _T_1939; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_1963 = _T_1934 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1490 = {{7'd0}, _T_1922}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_1965 = _T_1963 + _GEN_1490; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_13; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1493 = {{1{spriteYPositionReg_13[9]}},spriteYPositionReg_13}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_1991; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_13 = _T_1991[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2015 = {{1{inSpriteY_13[10]}},inSpriteY_13}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2033 = inSpriteX_13; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2041 = {{2'd0}, _T_2033}; // @[Mux.scala 80:57]
  wire [11:0] _T_2045 = {{1{inSpriteY_13[10]}},inSpriteY_13}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2053 = {{2'd0}, _T_2045}; // @[Mux.scala 80:57]
  wire  _T_2054 = $signed(inSpriteX_13) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2055 = $signed(inSpriteX_13) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2056 = _T_2054 & _T_2055; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2057 = $signed(_T_2015) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2058 = $signed(_T_2015) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2059 = _T_2057 & _T_2058; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2082 = _T_2053 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1499 = {{7'd0}, _T_2041}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2084 = _T_2082 + _GEN_1499; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_14; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1502 = {{1{spriteYPositionReg_14[9]}},spriteYPositionReg_14}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2110; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_14 = _T_2110[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2134 = {{1{inSpriteY_14[10]}},inSpriteY_14}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2152 = inSpriteX_14; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2160 = {{2'd0}, _T_2152}; // @[Mux.scala 80:57]
  wire [11:0] _T_2164 = {{1{inSpriteY_14[10]}},inSpriteY_14}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2172 = {{2'd0}, _T_2164}; // @[Mux.scala 80:57]
  wire  _T_2173 = $signed(inSpriteX_14) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2174 = $signed(inSpriteX_14) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2175 = _T_2173 & _T_2174; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2176 = $signed(_T_2134) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2177 = $signed(_T_2134) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2178 = _T_2176 & _T_2177; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2201 = _T_2172 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1508 = {{7'd0}, _T_2160}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2203 = _T_2201 + _GEN_1508; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_15; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1511 = {{1{spriteYPositionReg_15[9]}},spriteYPositionReg_15}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2229; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_15 = _T_2229[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2253 = {{1{inSpriteY_15[10]}},inSpriteY_15}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2271 = inSpriteX_15; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2279 = {{2'd0}, _T_2271}; // @[Mux.scala 80:57]
  wire [11:0] _T_2283 = {{1{inSpriteY_15[10]}},inSpriteY_15}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2291 = {{2'd0}, _T_2283}; // @[Mux.scala 80:57]
  wire  _T_2292 = $signed(inSpriteX_15) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2293 = $signed(inSpriteX_15) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2294 = _T_2292 & _T_2293; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2295 = $signed(_T_2253) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2296 = $signed(_T_2253) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2297 = _T_2295 & _T_2296; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2320 = _T_2291 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1517 = {{7'd0}, _T_2279}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2322 = _T_2320 + _GEN_1517; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_16; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1520 = {{1{spriteYPositionReg_16[9]}},spriteYPositionReg_16}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2348; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_16 = _T_2348[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2372 = {{1{inSpriteY_16[10]}},inSpriteY_16}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2390 = inSpriteX_16; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2398 = {{2'd0}, _T_2390}; // @[Mux.scala 80:57]
  wire [11:0] _T_2402 = {{1{inSpriteY_16[10]}},inSpriteY_16}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2410 = {{2'd0}, _T_2402}; // @[Mux.scala 80:57]
  wire  _T_2411 = $signed(inSpriteX_16) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2412 = $signed(inSpriteX_16) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2413 = _T_2411 & _T_2412; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2414 = $signed(_T_2372) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2415 = $signed(_T_2372) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2416 = _T_2414 & _T_2415; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2439 = _T_2410 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1526 = {{7'd0}, _T_2398}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2441 = _T_2439 + _GEN_1526; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_17; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1529 = {{1{spriteYPositionReg_17[9]}},spriteYPositionReg_17}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2467; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_17 = _T_2467[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2491 = {{1{inSpriteY_17[10]}},inSpriteY_17}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2509 = inSpriteX_17; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2517 = {{2'd0}, _T_2509}; // @[Mux.scala 80:57]
  wire [11:0] _T_2521 = {{1{inSpriteY_17[10]}},inSpriteY_17}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2529 = {{2'd0}, _T_2521}; // @[Mux.scala 80:57]
  wire  _T_2530 = $signed(inSpriteX_17) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2531 = $signed(inSpriteX_17) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2532 = _T_2530 & _T_2531; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2533 = $signed(_T_2491) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2534 = $signed(_T_2491) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2535 = _T_2533 & _T_2534; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2558 = _T_2529 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1535 = {{7'd0}, _T_2517}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2560 = _T_2558 + _GEN_1535; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_18; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1538 = {{1{spriteYPositionReg_18[9]}},spriteYPositionReg_18}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2586; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_18 = _T_2586[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2610 = {{1{inSpriteY_18[10]}},inSpriteY_18}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2628 = inSpriteX_18; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2636 = {{2'd0}, _T_2628}; // @[Mux.scala 80:57]
  wire [11:0] _T_2640 = {{1{inSpriteY_18[10]}},inSpriteY_18}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2648 = {{2'd0}, _T_2640}; // @[Mux.scala 80:57]
  wire  _T_2649 = $signed(inSpriteX_18) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2650 = $signed(inSpriteX_18) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2651 = _T_2649 & _T_2650; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2652 = $signed(_T_2610) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2653 = $signed(_T_2610) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2654 = _T_2652 & _T_2653; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2677 = _T_2648 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1544 = {{7'd0}, _T_2636}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2679 = _T_2677 + _GEN_1544; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_19; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1547 = {{1{spriteYPositionReg_19[9]}},spriteYPositionReg_19}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2705; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_19 = _T_2705[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2729 = {{1{inSpriteY_19[10]}},inSpriteY_19}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2747 = inSpriteX_19; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2755 = {{2'd0}, _T_2747}; // @[Mux.scala 80:57]
  wire [11:0] _T_2759 = {{1{inSpriteY_19[10]}},inSpriteY_19}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2767 = {{2'd0}, _T_2759}; // @[Mux.scala 80:57]
  wire  _T_2768 = $signed(inSpriteX_19) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2769 = $signed(inSpriteX_19) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2770 = _T_2768 & _T_2769; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2771 = $signed(_T_2729) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2772 = $signed(_T_2729) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2773 = _T_2771 & _T_2772; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2796 = _T_2767 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1553 = {{7'd0}, _T_2755}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2798 = _T_2796 + _GEN_1553; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_20; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1556 = {{1{spriteYPositionReg_20[9]}},spriteYPositionReg_20}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2824; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_20 = _T_2824[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2848 = {{1{inSpriteY_20[10]}},inSpriteY_20}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2866 = inSpriteX_20; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2874 = {{2'd0}, _T_2866}; // @[Mux.scala 80:57]
  wire [11:0] _T_2878 = {{1{inSpriteY_20[10]}},inSpriteY_20}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_2886 = {{2'd0}, _T_2878}; // @[Mux.scala 80:57]
  wire  _T_2887 = $signed(inSpriteX_20) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_2888 = $signed(inSpriteX_20) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_2889 = _T_2887 & _T_2888; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_2890 = $signed(_T_2848) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_2891 = $signed(_T_2848) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_2892 = _T_2890 & _T_2891; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_2915 = _T_2886 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1562 = {{7'd0}, _T_2874}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_2917 = _T_2915 + _GEN_1562; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_21; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1565 = {{1{spriteYPositionReg_21[9]}},spriteYPositionReg_21}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_2943; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_21 = _T_2943[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_2967 = {{1{inSpriteY_21[10]}},inSpriteY_21}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_2985 = inSpriteX_21; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_2993 = {{2'd0}, _T_2985}; // @[Mux.scala 80:57]
  wire [11:0] _T_2997 = {{1{inSpriteY_21[10]}},inSpriteY_21}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3005 = {{2'd0}, _T_2997}; // @[Mux.scala 80:57]
  wire  _T_3006 = $signed(inSpriteX_21) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3007 = $signed(inSpriteX_21) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3008 = _T_3006 & _T_3007; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3009 = $signed(_T_2967) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3010 = $signed(_T_2967) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3011 = _T_3009 & _T_3010; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3034 = _T_3005 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1571 = {{7'd0}, _T_2993}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3036 = _T_3034 + _GEN_1571; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_22; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1574 = {{1{spriteYPositionReg_22[9]}},spriteYPositionReg_22}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3062; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_22 = _T_3062[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3086 = {{1{inSpriteY_22[10]}},inSpriteY_22}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3104 = inSpriteX_22; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3112 = {{2'd0}, _T_3104}; // @[Mux.scala 80:57]
  wire [11:0] _T_3116 = {{1{inSpriteY_22[10]}},inSpriteY_22}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3124 = {{2'd0}, _T_3116}; // @[Mux.scala 80:57]
  wire  _T_3125 = $signed(inSpriteX_22) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3126 = $signed(inSpriteX_22) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3127 = _T_3125 & _T_3126; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3128 = $signed(_T_3086) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3129 = $signed(_T_3086) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3130 = _T_3128 & _T_3129; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3153 = _T_3124 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1580 = {{7'd0}, _T_3112}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3155 = _T_3153 + _GEN_1580; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_23; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1583 = {{1{spriteYPositionReg_23[9]}},spriteYPositionReg_23}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3181; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_23 = _T_3181[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3205 = {{1{inSpriteY_23[10]}},inSpriteY_23}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3223 = inSpriteX_23; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3231 = {{2'd0}, _T_3223}; // @[Mux.scala 80:57]
  wire [11:0] _T_3235 = {{1{inSpriteY_23[10]}},inSpriteY_23}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3243 = {{2'd0}, _T_3235}; // @[Mux.scala 80:57]
  wire  _T_3244 = $signed(inSpriteX_23) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3245 = $signed(inSpriteX_23) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3246 = _T_3244 & _T_3245; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3247 = $signed(_T_3205) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3248 = $signed(_T_3205) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3249 = _T_3247 & _T_3248; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3272 = _T_3243 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1589 = {{7'd0}, _T_3231}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3274 = _T_3272 + _GEN_1589; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_24; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1592 = {{1{spriteYPositionReg_24[9]}},spriteYPositionReg_24}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3300; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_24 = _T_3300[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3324 = {{1{inSpriteY_24[10]}},inSpriteY_24}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3342 = inSpriteX_24; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3350 = {{2'd0}, _T_3342}; // @[Mux.scala 80:57]
  wire [11:0] _T_3354 = {{1{inSpriteY_24[10]}},inSpriteY_24}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3362 = {{2'd0}, _T_3354}; // @[Mux.scala 80:57]
  wire  _T_3363 = $signed(inSpriteX_24) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3364 = $signed(inSpriteX_24) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3365 = _T_3363 & _T_3364; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3366 = $signed(_T_3324) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3367 = $signed(_T_3324) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3368 = _T_3366 & _T_3367; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3391 = _T_3362 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1598 = {{7'd0}, _T_3350}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3393 = _T_3391 + _GEN_1598; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_25; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1601 = {{1{spriteYPositionReg_25[9]}},spriteYPositionReg_25}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3419; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_25 = _T_3419[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3443 = {{1{inSpriteY_25[10]}},inSpriteY_25}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3461 = inSpriteX_25; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3469 = {{2'd0}, _T_3461}; // @[Mux.scala 80:57]
  wire [11:0] _T_3473 = {{1{inSpriteY_25[10]}},inSpriteY_25}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3481 = {{2'd0}, _T_3473}; // @[Mux.scala 80:57]
  wire  _T_3482 = $signed(inSpriteX_25) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3483 = $signed(inSpriteX_25) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3484 = _T_3482 & _T_3483; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3485 = $signed(_T_3443) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3486 = $signed(_T_3443) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3487 = _T_3485 & _T_3486; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3510 = _T_3481 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1607 = {{7'd0}, _T_3469}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3512 = _T_3510 + _GEN_1607; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_26; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1610 = {{1{spriteYPositionReg_26[9]}},spriteYPositionReg_26}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3538; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_26 = _T_3538[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3562 = {{1{inSpriteY_26[10]}},inSpriteY_26}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3580 = inSpriteX_26; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3588 = {{2'd0}, _T_3580}; // @[Mux.scala 80:57]
  wire [11:0] _T_3592 = {{1{inSpriteY_26[10]}},inSpriteY_26}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3600 = {{2'd0}, _T_3592}; // @[Mux.scala 80:57]
  wire  _T_3601 = $signed(inSpriteX_26) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3602 = $signed(inSpriteX_26) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3603 = _T_3601 & _T_3602; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3604 = $signed(_T_3562) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3605 = $signed(_T_3562) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3606 = _T_3604 & _T_3605; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3629 = _T_3600 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1616 = {{7'd0}, _T_3588}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3631 = _T_3629 + _GEN_1616; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_27; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1619 = {{1{spriteYPositionReg_27[9]}},spriteYPositionReg_27}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3657; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_27 = _T_3657[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3681 = {{1{inSpriteY_27[10]}},inSpriteY_27}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3699 = inSpriteX_27; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3707 = {{2'd0}, _T_3699}; // @[Mux.scala 80:57]
  wire [11:0] _T_3711 = {{1{inSpriteY_27[10]}},inSpriteY_27}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3719 = {{2'd0}, _T_3711}; // @[Mux.scala 80:57]
  wire  _T_3720 = $signed(inSpriteX_27) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3721 = $signed(inSpriteX_27) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3722 = _T_3720 & _T_3721; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3723 = $signed(_T_3681) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3724 = $signed(_T_3681) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3725 = _T_3723 & _T_3724; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3748 = _T_3719 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1625 = {{7'd0}, _T_3707}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3750 = _T_3748 + _GEN_1625; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_28; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1628 = {{1{spriteYPositionReg_28[9]}},spriteYPositionReg_28}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3776; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_28 = _T_3776[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3800 = {{1{inSpriteY_28[10]}},inSpriteY_28}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3818 = inSpriteX_28; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3826 = {{2'd0}, _T_3818}; // @[Mux.scala 80:57]
  wire [11:0] _T_3830 = {{1{inSpriteY_28[10]}},inSpriteY_28}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3838 = {{2'd0}, _T_3830}; // @[Mux.scala 80:57]
  wire  _T_3839 = $signed(inSpriteX_28) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3840 = $signed(inSpriteX_28) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3841 = _T_3839 & _T_3840; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3842 = $signed(_T_3800) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3843 = $signed(_T_3800) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3844 = _T_3842 & _T_3843; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3867 = _T_3838 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1634 = {{7'd0}, _T_3826}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3869 = _T_3867 + _GEN_1634; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_29; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1637 = {{1{spriteYPositionReg_29[9]}},spriteYPositionReg_29}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_3895; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_29 = _T_3895[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_3919 = {{1{inSpriteY_29[10]}},inSpriteY_29}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_3937 = inSpriteX_29; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_3945 = {{2'd0}, _T_3937}; // @[Mux.scala 80:57]
  wire [11:0] _T_3949 = {{1{inSpriteY_29[10]}},inSpriteY_29}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_3957 = {{2'd0}, _T_3949}; // @[Mux.scala 80:57]
  wire  _T_3958 = $signed(inSpriteX_29) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_3959 = $signed(inSpriteX_29) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_3960 = _T_3958 & _T_3959; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_3961 = $signed(_T_3919) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_3962 = $signed(_T_3919) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_3963 = _T_3961 & _T_3962; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_3986 = _T_3957 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1643 = {{7'd0}, _T_3945}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_3988 = _T_3986 + _GEN_1643; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_30; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1646 = {{1{spriteYPositionReg_30[9]}},spriteYPositionReg_30}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4014; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_30 = _T_4014[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4038 = {{1{inSpriteY_30[10]}},inSpriteY_30}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4056 = inSpriteX_30; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4064 = {{2'd0}, _T_4056}; // @[Mux.scala 80:57]
  wire [11:0] _T_4068 = {{1{inSpriteY_30[10]}},inSpriteY_30}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4076 = {{2'd0}, _T_4068}; // @[Mux.scala 80:57]
  wire  _T_4077 = $signed(inSpriteX_30) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4078 = $signed(inSpriteX_30) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4079 = _T_4077 & _T_4078; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4080 = $signed(_T_4038) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4081 = $signed(_T_4038) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4082 = _T_4080 & _T_4081; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4105 = _T_4076 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1652 = {{7'd0}, _T_4064}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4107 = _T_4105 + _GEN_1652; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_31; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1655 = {{1{spriteYPositionReg_31[9]}},spriteYPositionReg_31}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4133; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_31 = _T_4133[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4157 = {{1{inSpriteY_31[10]}},inSpriteY_31}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4175 = inSpriteX_31; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4183 = {{2'd0}, _T_4175}; // @[Mux.scala 80:57]
  wire [11:0] _T_4187 = {{1{inSpriteY_31[10]}},inSpriteY_31}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4195 = {{2'd0}, _T_4187}; // @[Mux.scala 80:57]
  wire  _T_4196 = $signed(inSpriteX_31) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4197 = $signed(inSpriteX_31) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4198 = _T_4196 & _T_4197; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4199 = $signed(_T_4157) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4200 = $signed(_T_4157) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4201 = _T_4199 & _T_4200; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4224 = _T_4195 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1661 = {{7'd0}, _T_4183}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4226 = _T_4224 + _GEN_1661; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_32; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1664 = {{1{spriteYPositionReg_32[9]}},spriteYPositionReg_32}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4252; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_32 = _T_4252[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4276 = {{1{inSpriteY_32[10]}},inSpriteY_32}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4294 = inSpriteX_32; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4302 = {{2'd0}, _T_4294}; // @[Mux.scala 80:57]
  wire [11:0] _T_4306 = {{1{inSpriteY_32[10]}},inSpriteY_32}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4314 = {{2'd0}, _T_4306}; // @[Mux.scala 80:57]
  wire  _T_4315 = $signed(inSpriteX_32) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4316 = $signed(inSpriteX_32) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4317 = _T_4315 & _T_4316; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4318 = $signed(_T_4276) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4319 = $signed(_T_4276) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4320 = _T_4318 & _T_4319; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4343 = _T_4314 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1670 = {{7'd0}, _T_4302}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4345 = _T_4343 + _GEN_1670; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_33; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1673 = {{1{spriteYPositionReg_33[9]}},spriteYPositionReg_33}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4371; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_33 = _T_4371[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4395 = {{1{inSpriteY_33[10]}},inSpriteY_33}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4413 = inSpriteX_33; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4421 = {{2'd0}, _T_4413}; // @[Mux.scala 80:57]
  wire [11:0] _T_4425 = {{1{inSpriteY_33[10]}},inSpriteY_33}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4433 = {{2'd0}, _T_4425}; // @[Mux.scala 80:57]
  wire  _T_4434 = $signed(inSpriteX_33) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4435 = $signed(inSpriteX_33) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4436 = _T_4434 & _T_4435; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4437 = $signed(_T_4395) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4438 = $signed(_T_4395) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4439 = _T_4437 & _T_4438; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4462 = _T_4433 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1679 = {{7'd0}, _T_4421}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4464 = _T_4462 + _GEN_1679; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_34; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1682 = {{1{spriteYPositionReg_34[9]}},spriteYPositionReg_34}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4490; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_34 = _T_4490[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4514 = {{1{inSpriteY_34[10]}},inSpriteY_34}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4532 = inSpriteX_34; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4540 = {{2'd0}, _T_4532}; // @[Mux.scala 80:57]
  wire [11:0] _T_4544 = {{1{inSpriteY_34[10]}},inSpriteY_34}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4552 = {{2'd0}, _T_4544}; // @[Mux.scala 80:57]
  wire  _T_4553 = $signed(inSpriteX_34) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4554 = $signed(inSpriteX_34) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4555 = _T_4553 & _T_4554; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4556 = $signed(_T_4514) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4557 = $signed(_T_4514) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4558 = _T_4556 & _T_4557; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4581 = _T_4552 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1688 = {{7'd0}, _T_4540}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4583 = _T_4581 + _GEN_1688; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_35; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1691 = {{1{spriteYPositionReg_35[9]}},spriteYPositionReg_35}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4609; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_35 = _T_4609[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4633 = {{1{inSpriteY_35[10]}},inSpriteY_35}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4651 = inSpriteX_35; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4659 = {{2'd0}, _T_4651}; // @[Mux.scala 80:57]
  wire [11:0] _T_4663 = {{1{inSpriteY_35[10]}},inSpriteY_35}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4671 = {{2'd0}, _T_4663}; // @[Mux.scala 80:57]
  wire  _T_4672 = $signed(inSpriteX_35) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4673 = $signed(inSpriteX_35) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4674 = _T_4672 & _T_4673; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4675 = $signed(_T_4633) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4676 = $signed(_T_4633) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4677 = _T_4675 & _T_4676; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4700 = _T_4671 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1697 = {{7'd0}, _T_4659}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4702 = _T_4700 + _GEN_1697; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_36; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1700 = {{1{spriteYPositionReg_36[9]}},spriteYPositionReg_36}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4728; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_36 = _T_4728[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4752 = {{1{inSpriteY_36[10]}},inSpriteY_36}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4770 = inSpriteX_36; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4778 = {{2'd0}, _T_4770}; // @[Mux.scala 80:57]
  wire [11:0] _T_4782 = {{1{inSpriteY_36[10]}},inSpriteY_36}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4790 = {{2'd0}, _T_4782}; // @[Mux.scala 80:57]
  wire  _T_4791 = $signed(inSpriteX_36) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4792 = $signed(inSpriteX_36) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4793 = _T_4791 & _T_4792; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4794 = $signed(_T_4752) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4795 = $signed(_T_4752) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4796 = _T_4794 & _T_4795; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4819 = _T_4790 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1706 = {{7'd0}, _T_4778}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4821 = _T_4819 + _GEN_1706; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_37; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1709 = {{1{spriteYPositionReg_37[9]}},spriteYPositionReg_37}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4847; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_37 = _T_4847[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4871 = {{1{inSpriteY_37[10]}},inSpriteY_37}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_4889 = inSpriteX_37; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_4897 = {{2'd0}, _T_4889}; // @[Mux.scala 80:57]
  wire [11:0] _T_4901 = {{1{inSpriteY_37[10]}},inSpriteY_37}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_4909 = {{2'd0}, _T_4901}; // @[Mux.scala 80:57]
  wire  _T_4910 = $signed(inSpriteX_37) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_4911 = $signed(inSpriteX_37) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_4912 = _T_4910 & _T_4911; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_4913 = $signed(_T_4871) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_4914 = $signed(_T_4871) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_4915 = _T_4913 & _T_4914; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_4938 = _T_4909 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1715 = {{7'd0}, _T_4897}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_4940 = _T_4938 + _GEN_1715; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_38; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1718 = {{1{spriteYPositionReg_38[9]}},spriteYPositionReg_38}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_4966; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_38 = _T_4966[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_4990 = {{1{inSpriteY_38[10]}},inSpriteY_38}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5008 = inSpriteX_38; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5016 = {{2'd0}, _T_5008}; // @[Mux.scala 80:57]
  wire [11:0] _T_5020 = {{1{inSpriteY_38[10]}},inSpriteY_38}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5028 = {{2'd0}, _T_5020}; // @[Mux.scala 80:57]
  wire  _T_5029 = $signed(inSpriteX_38) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5030 = $signed(inSpriteX_38) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5031 = _T_5029 & _T_5030; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5032 = $signed(_T_4990) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5033 = $signed(_T_4990) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5034 = _T_5032 & _T_5033; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5057 = _T_5028 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1724 = {{7'd0}, _T_5016}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5059 = _T_5057 + _GEN_1724; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_39; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1727 = {{1{spriteYPositionReg_39[9]}},spriteYPositionReg_39}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5085; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_39 = _T_5085[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5109 = {{1{inSpriteY_39[10]}},inSpriteY_39}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5127 = inSpriteX_39; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5135 = {{2'd0}, _T_5127}; // @[Mux.scala 80:57]
  wire [11:0] _T_5139 = {{1{inSpriteY_39[10]}},inSpriteY_39}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5147 = {{2'd0}, _T_5139}; // @[Mux.scala 80:57]
  wire  _T_5148 = $signed(inSpriteX_39) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5149 = $signed(inSpriteX_39) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5150 = _T_5148 & _T_5149; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5151 = $signed(_T_5109) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5152 = $signed(_T_5109) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5153 = _T_5151 & _T_5152; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5176 = _T_5147 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1733 = {{7'd0}, _T_5135}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5178 = _T_5176 + _GEN_1733; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_40; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1736 = {{1{spriteYPositionReg_40[9]}},spriteYPositionReg_40}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5204; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_40 = _T_5204[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5228 = {{1{inSpriteY_40[10]}},inSpriteY_40}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5246 = inSpriteX_40; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5254 = {{2'd0}, _T_5246}; // @[Mux.scala 80:57]
  wire [11:0] _T_5258 = {{1{inSpriteY_40[10]}},inSpriteY_40}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5266 = {{2'd0}, _T_5258}; // @[Mux.scala 80:57]
  wire  _T_5267 = $signed(inSpriteX_40) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5268 = $signed(inSpriteX_40) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5269 = _T_5267 & _T_5268; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5270 = $signed(_T_5228) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5271 = $signed(_T_5228) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5272 = _T_5270 & _T_5271; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5295 = _T_5266 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1742 = {{7'd0}, _T_5254}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5297 = _T_5295 + _GEN_1742; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_41; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1745 = {{1{spriteYPositionReg_41[9]}},spriteYPositionReg_41}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5323; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_41 = _T_5323[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5347 = {{1{inSpriteY_41[10]}},inSpriteY_41}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5365 = inSpriteX_41; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5373 = {{2'd0}, _T_5365}; // @[Mux.scala 80:57]
  wire [11:0] _T_5377 = {{1{inSpriteY_41[10]}},inSpriteY_41}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5385 = {{2'd0}, _T_5377}; // @[Mux.scala 80:57]
  wire  _T_5386 = $signed(inSpriteX_41) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5387 = $signed(inSpriteX_41) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5388 = _T_5386 & _T_5387; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5389 = $signed(_T_5347) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5390 = $signed(_T_5347) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5391 = _T_5389 & _T_5390; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5414 = _T_5385 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1751 = {{7'd0}, _T_5373}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5416 = _T_5414 + _GEN_1751; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_42; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1754 = {{1{spriteYPositionReg_42[9]}},spriteYPositionReg_42}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5442; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_42 = _T_5442[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5466 = {{1{inSpriteY_42[10]}},inSpriteY_42}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5484 = inSpriteX_42; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5492 = {{2'd0}, _T_5484}; // @[Mux.scala 80:57]
  wire [11:0] _T_5496 = {{1{inSpriteY_42[10]}},inSpriteY_42}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5504 = {{2'd0}, _T_5496}; // @[Mux.scala 80:57]
  wire  _T_5505 = $signed(inSpriteX_42) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5506 = $signed(inSpriteX_42) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5507 = _T_5505 & _T_5506; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5508 = $signed(_T_5466) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5509 = $signed(_T_5466) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5510 = _T_5508 & _T_5509; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5533 = _T_5504 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1760 = {{7'd0}, _T_5492}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5535 = _T_5533 + _GEN_1760; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_43; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1763 = {{1{spriteYPositionReg_43[9]}},spriteYPositionReg_43}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5561; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_43 = _T_5561[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5585 = {{1{inSpriteY_43[10]}},inSpriteY_43}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5603 = inSpriteX_43; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5611 = {{2'd0}, _T_5603}; // @[Mux.scala 80:57]
  wire [11:0] _T_5615 = {{1{inSpriteY_43[10]}},inSpriteY_43}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5623 = {{2'd0}, _T_5615}; // @[Mux.scala 80:57]
  wire  _T_5624 = $signed(inSpriteX_43) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5625 = $signed(inSpriteX_43) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5626 = _T_5624 & _T_5625; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5627 = $signed(_T_5585) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5628 = $signed(_T_5585) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5629 = _T_5627 & _T_5628; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5652 = _T_5623 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1769 = {{7'd0}, _T_5611}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5654 = _T_5652 + _GEN_1769; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_44; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1772 = {{1{spriteYPositionReg_44[9]}},spriteYPositionReg_44}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5680; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_44 = _T_5680[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5704 = {{1{inSpriteY_44[10]}},inSpriteY_44}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5722 = inSpriteX_44; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5730 = {{2'd0}, _T_5722}; // @[Mux.scala 80:57]
  wire [11:0] _T_5734 = {{1{inSpriteY_44[10]}},inSpriteY_44}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5742 = {{2'd0}, _T_5734}; // @[Mux.scala 80:57]
  wire  _T_5743 = $signed(inSpriteX_44) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5744 = $signed(inSpriteX_44) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5745 = _T_5743 & _T_5744; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5746 = $signed(_T_5704) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5747 = $signed(_T_5704) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5748 = _T_5746 & _T_5747; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5771 = _T_5742 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1778 = {{7'd0}, _T_5730}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5773 = _T_5771 + _GEN_1778; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_45; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1781 = {{1{spriteYPositionReg_45[9]}},spriteYPositionReg_45}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5799; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_45 = _T_5799[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5823 = {{1{inSpriteY_45[10]}},inSpriteY_45}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5841 = inSpriteX_45; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5849 = {{2'd0}, _T_5841}; // @[Mux.scala 80:57]
  wire [11:0] _T_5853 = {{1{inSpriteY_45[10]}},inSpriteY_45}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5861 = {{2'd0}, _T_5853}; // @[Mux.scala 80:57]
  wire  _T_5862 = $signed(inSpriteX_45) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5863 = $signed(inSpriteX_45) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5864 = _T_5862 & _T_5863; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5865 = $signed(_T_5823) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5866 = $signed(_T_5823) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5867 = _T_5865 & _T_5866; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_5890 = _T_5861 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1787 = {{7'd0}, _T_5849}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_5892 = _T_5890 + _GEN_1787; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_46; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1790 = {{1{spriteYPositionReg_46[9]}},spriteYPositionReg_46}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_5918; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_46 = _T_5918[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_5942 = {{1{inSpriteY_46[10]}},inSpriteY_46}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_5960 = inSpriteX_46; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_5968 = {{2'd0}, _T_5960}; // @[Mux.scala 80:57]
  wire [11:0] _T_5972 = {{1{inSpriteY_46[10]}},inSpriteY_46}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_5980 = {{2'd0}, _T_5972}; // @[Mux.scala 80:57]
  wire  _T_5981 = $signed(inSpriteX_46) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_5982 = $signed(inSpriteX_46) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_5983 = _T_5981 & _T_5982; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_5984 = $signed(_T_5942) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_5985 = $signed(_T_5942) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_5986 = _T_5984 & _T_5985; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6009 = _T_5980 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1796 = {{7'd0}, _T_5968}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6011 = _T_6009 + _GEN_1796; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_47; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1799 = {{1{spriteYPositionReg_47[9]}},spriteYPositionReg_47}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6037; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_47 = _T_6037[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6061 = {{1{inSpriteY_47[10]}},inSpriteY_47}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6079 = inSpriteX_47; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6087 = {{2'd0}, _T_6079}; // @[Mux.scala 80:57]
  wire [11:0] _T_6091 = {{1{inSpriteY_47[10]}},inSpriteY_47}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6099 = {{2'd0}, _T_6091}; // @[Mux.scala 80:57]
  wire  _T_6100 = $signed(inSpriteX_47) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6101 = $signed(inSpriteX_47) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6102 = _T_6100 & _T_6101; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6103 = $signed(_T_6061) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6104 = $signed(_T_6061) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6105 = _T_6103 & _T_6104; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6128 = _T_6099 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1805 = {{7'd0}, _T_6087}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6130 = _T_6128 + _GEN_1805; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_48; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1808 = {{1{spriteYPositionReg_48[9]}},spriteYPositionReg_48}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6156; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_48 = _T_6156[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6180 = {{1{inSpriteY_48[10]}},inSpriteY_48}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6198 = inSpriteX_48; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6206 = {{2'd0}, _T_6198}; // @[Mux.scala 80:57]
  wire [11:0] _T_6210 = {{1{inSpriteY_48[10]}},inSpriteY_48}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6218 = {{2'd0}, _T_6210}; // @[Mux.scala 80:57]
  wire  _T_6219 = $signed(inSpriteX_48) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6220 = $signed(inSpriteX_48) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6221 = _T_6219 & _T_6220; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6222 = $signed(_T_6180) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6223 = $signed(_T_6180) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6224 = _T_6222 & _T_6223; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6247 = _T_6218 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1814 = {{7'd0}, _T_6206}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6249 = _T_6247 + _GEN_1814; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_49; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1817 = {{1{spriteYPositionReg_49[9]}},spriteYPositionReg_49}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6275; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_49 = _T_6275[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6299 = {{1{inSpriteY_49[10]}},inSpriteY_49}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6317 = inSpriteX_49; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6325 = {{2'd0}, _T_6317}; // @[Mux.scala 80:57]
  wire [11:0] _T_6329 = {{1{inSpriteY_49[10]}},inSpriteY_49}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6337 = {{2'd0}, _T_6329}; // @[Mux.scala 80:57]
  wire  _T_6338 = $signed(inSpriteX_49) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6339 = $signed(inSpriteX_49) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6340 = _T_6338 & _T_6339; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6341 = $signed(_T_6299) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6342 = $signed(_T_6299) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6343 = _T_6341 & _T_6342; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6366 = _T_6337 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1823 = {{7'd0}, _T_6325}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6368 = _T_6366 + _GEN_1823; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_50; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1826 = {{1{spriteYPositionReg_50[9]}},spriteYPositionReg_50}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6394; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_50 = _T_6394[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6418 = {{1{inSpriteY_50[10]}},inSpriteY_50}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6436 = inSpriteX_50; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6444 = {{2'd0}, _T_6436}; // @[Mux.scala 80:57]
  wire [11:0] _T_6448 = {{1{inSpriteY_50[10]}},inSpriteY_50}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6456 = {{2'd0}, _T_6448}; // @[Mux.scala 80:57]
  wire  _T_6457 = $signed(inSpriteX_50) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6458 = $signed(inSpriteX_50) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6459 = _T_6457 & _T_6458; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6460 = $signed(_T_6418) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6461 = $signed(_T_6418) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6462 = _T_6460 & _T_6461; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6485 = _T_6456 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1832 = {{7'd0}, _T_6444}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6487 = _T_6485 + _GEN_1832; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_51; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1835 = {{1{spriteYPositionReg_51[9]}},spriteYPositionReg_51}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6513; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_51 = _T_6513[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6537 = {{1{inSpriteY_51[10]}},inSpriteY_51}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6555 = inSpriteX_51; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6563 = {{2'd0}, _T_6555}; // @[Mux.scala 80:57]
  wire [11:0] _T_6567 = {{1{inSpriteY_51[10]}},inSpriteY_51}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6575 = {{2'd0}, _T_6567}; // @[Mux.scala 80:57]
  wire  _T_6576 = $signed(inSpriteX_51) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6577 = $signed(inSpriteX_51) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6578 = _T_6576 & _T_6577; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6579 = $signed(_T_6537) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6580 = $signed(_T_6537) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6581 = _T_6579 & _T_6580; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6604 = _T_6575 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1841 = {{7'd0}, _T_6563}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6606 = _T_6604 + _GEN_1841; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_52; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1844 = {{1{spriteYPositionReg_52[9]}},spriteYPositionReg_52}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6632; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_52 = _T_6632[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6656 = {{1{inSpriteY_52[10]}},inSpriteY_52}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6674 = inSpriteX_52; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6682 = {{2'd0}, _T_6674}; // @[Mux.scala 80:57]
  wire [11:0] _T_6686 = {{1{inSpriteY_52[10]}},inSpriteY_52}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6694 = {{2'd0}, _T_6686}; // @[Mux.scala 80:57]
  wire  _T_6695 = $signed(inSpriteX_52) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6696 = $signed(inSpriteX_52) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6697 = _T_6695 & _T_6696; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6698 = $signed(_T_6656) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6699 = $signed(_T_6656) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6700 = _T_6698 & _T_6699; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6723 = _T_6694 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1850 = {{7'd0}, _T_6682}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6725 = _T_6723 + _GEN_1850; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_53; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1853 = {{1{spriteYPositionReg_53[9]}},spriteYPositionReg_53}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6751; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_53 = _T_6751[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6775 = {{1{inSpriteY_53[10]}},inSpriteY_53}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6793 = inSpriteX_53; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6801 = {{2'd0}, _T_6793}; // @[Mux.scala 80:57]
  wire [11:0] _T_6805 = {{1{inSpriteY_53[10]}},inSpriteY_53}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6813 = {{2'd0}, _T_6805}; // @[Mux.scala 80:57]
  wire  _T_6814 = $signed(inSpriteX_53) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6815 = $signed(inSpriteX_53) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6816 = _T_6814 & _T_6815; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6817 = $signed(_T_6775) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6818 = $signed(_T_6775) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6819 = _T_6817 & _T_6818; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6842 = _T_6813 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1859 = {{7'd0}, _T_6801}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6844 = _T_6842 + _GEN_1859; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_54; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1862 = {{1{spriteYPositionReg_54[9]}},spriteYPositionReg_54}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6870; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_54 = _T_6870[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_6894 = {{1{inSpriteY_54[10]}},inSpriteY_54}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_6912 = inSpriteX_54; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_6920 = {{2'd0}, _T_6912}; // @[Mux.scala 80:57]
  wire [11:0] _T_6924 = {{1{inSpriteY_54[10]}},inSpriteY_54}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_6932 = {{2'd0}, _T_6924}; // @[Mux.scala 80:57]
  wire  _T_6933 = $signed(inSpriteX_54) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_6934 = $signed(inSpriteX_54) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_6935 = _T_6933 & _T_6934; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_6936 = $signed(_T_6894) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_6937 = $signed(_T_6894) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_6938 = _T_6936 & _T_6937; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_6961 = _T_6932 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1868 = {{7'd0}, _T_6920}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_6963 = _T_6961 + _GEN_1868; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_55; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1871 = {{1{spriteYPositionReg_55[9]}},spriteYPositionReg_55}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_6989; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_55 = _T_6989[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7013 = {{1{inSpriteY_55[10]}},inSpriteY_55}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7031 = inSpriteX_55; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7039 = {{2'd0}, _T_7031}; // @[Mux.scala 80:57]
  wire [11:0] _T_7043 = {{1{inSpriteY_55[10]}},inSpriteY_55}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7051 = {{2'd0}, _T_7043}; // @[Mux.scala 80:57]
  wire  _T_7052 = $signed(inSpriteX_55) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7053 = $signed(inSpriteX_55) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7054 = _T_7052 & _T_7053; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7055 = $signed(_T_7013) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7056 = $signed(_T_7013) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7057 = _T_7055 & _T_7056; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7080 = _T_7051 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1877 = {{7'd0}, _T_7039}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7082 = _T_7080 + _GEN_1877; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_56; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1880 = {{1{spriteYPositionReg_56[9]}},spriteYPositionReg_56}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7108; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_56 = _T_7108[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7132 = {{1{inSpriteY_56[10]}},inSpriteY_56}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7150 = inSpriteX_56; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7158 = {{2'd0}, _T_7150}; // @[Mux.scala 80:57]
  wire [11:0] _T_7162 = {{1{inSpriteY_56[10]}},inSpriteY_56}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7170 = {{2'd0}, _T_7162}; // @[Mux.scala 80:57]
  wire  _T_7171 = $signed(inSpriteX_56) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7172 = $signed(inSpriteX_56) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7173 = _T_7171 & _T_7172; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7174 = $signed(_T_7132) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7175 = $signed(_T_7132) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7176 = _T_7174 & _T_7175; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7199 = _T_7170 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1886 = {{7'd0}, _T_7158}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7201 = _T_7199 + _GEN_1886; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_57; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1889 = {{1{spriteYPositionReg_57[9]}},spriteYPositionReg_57}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7227; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_57 = _T_7227[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7251 = {{1{inSpriteY_57[10]}},inSpriteY_57}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7269 = inSpriteX_57; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7277 = {{2'd0}, _T_7269}; // @[Mux.scala 80:57]
  wire [11:0] _T_7281 = {{1{inSpriteY_57[10]}},inSpriteY_57}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7289 = {{2'd0}, _T_7281}; // @[Mux.scala 80:57]
  wire  _T_7290 = $signed(inSpriteX_57) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7291 = $signed(inSpriteX_57) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7292 = _T_7290 & _T_7291; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7293 = $signed(_T_7251) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7294 = $signed(_T_7251) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7295 = _T_7293 & _T_7294; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7318 = _T_7289 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1895 = {{7'd0}, _T_7277}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7320 = _T_7318 + _GEN_1895; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_58; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1898 = {{1{spriteYPositionReg_58[9]}},spriteYPositionReg_58}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7346; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_58 = _T_7346[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7370 = {{1{inSpriteY_58[10]}},inSpriteY_58}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7388 = inSpriteX_58; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7396 = {{2'd0}, _T_7388}; // @[Mux.scala 80:57]
  wire [11:0] _T_7400 = {{1{inSpriteY_58[10]}},inSpriteY_58}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7408 = {{2'd0}, _T_7400}; // @[Mux.scala 80:57]
  wire  _T_7409 = $signed(inSpriteX_58) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7410 = $signed(inSpriteX_58) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7411 = _T_7409 & _T_7410; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7412 = $signed(_T_7370) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7413 = $signed(_T_7370) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7414 = _T_7412 & _T_7413; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7437 = _T_7408 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1904 = {{7'd0}, _T_7396}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7439 = _T_7437 + _GEN_1904; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_59; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1907 = {{1{spriteYPositionReg_59[9]}},spriteYPositionReg_59}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7465; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_59 = _T_7465[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7489 = {{1{inSpriteY_59[10]}},inSpriteY_59}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7507 = inSpriteX_59; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7515 = {{2'd0}, _T_7507}; // @[Mux.scala 80:57]
  wire [11:0] _T_7519 = {{1{inSpriteY_59[10]}},inSpriteY_59}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7527 = {{2'd0}, _T_7519}; // @[Mux.scala 80:57]
  wire  _T_7528 = $signed(inSpriteX_59) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7529 = $signed(inSpriteX_59) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7530 = _T_7528 & _T_7529; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7531 = $signed(_T_7489) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7532 = $signed(_T_7489) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7533 = _T_7531 & _T_7532; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7556 = _T_7527 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1913 = {{7'd0}, _T_7515}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7558 = _T_7556 + _GEN_1913; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_60; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1916 = {{1{spriteYPositionReg_60[9]}},spriteYPositionReg_60}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7584; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_60 = _T_7584[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7608 = {{1{inSpriteY_60[10]}},inSpriteY_60}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7626 = inSpriteX_60; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7634 = {{2'd0}, _T_7626}; // @[Mux.scala 80:57]
  wire [11:0] _T_7638 = {{1{inSpriteY_60[10]}},inSpriteY_60}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7646 = {{2'd0}, _T_7638}; // @[Mux.scala 80:57]
  wire  _T_7647 = $signed(inSpriteX_60) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7648 = $signed(inSpriteX_60) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7649 = _T_7647 & _T_7648; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7650 = $signed(_T_7608) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7651 = $signed(_T_7608) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7652 = _T_7650 & _T_7651; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7675 = _T_7646 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1922 = {{7'd0}, _T_7634}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7677 = _T_7675 + _GEN_1922; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_61; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1925 = {{1{spriteYPositionReg_61[9]}},spriteYPositionReg_61}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7703; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_61 = _T_7703[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7727 = {{1{inSpriteY_61[10]}},inSpriteY_61}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7745 = inSpriteX_61; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7753 = {{2'd0}, _T_7745}; // @[Mux.scala 80:57]
  wire [11:0] _T_7757 = {{1{inSpriteY_61[10]}},inSpriteY_61}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7765 = {{2'd0}, _T_7757}; // @[Mux.scala 80:57]
  wire  _T_7766 = $signed(inSpriteX_61) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7767 = $signed(inSpriteX_61) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7768 = _T_7766 & _T_7767; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7769 = $signed(_T_7727) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7770 = $signed(_T_7727) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7771 = _T_7769 & _T_7770; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7794 = _T_7765 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1931 = {{7'd0}, _T_7753}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7796 = _T_7794 + _GEN_1931; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_62; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1934 = {{1{spriteYPositionReg_62[9]}},spriteYPositionReg_62}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7822; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_62 = _T_7822[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7846 = {{1{inSpriteY_62[10]}},inSpriteY_62}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7864 = inSpriteX_62; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7872 = {{2'd0}, _T_7864}; // @[Mux.scala 80:57]
  wire [11:0] _T_7876 = {{1{inSpriteY_62[10]}},inSpriteY_62}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_7884 = {{2'd0}, _T_7876}; // @[Mux.scala 80:57]
  wire  _T_7885 = $signed(inSpriteX_62) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_7886 = $signed(inSpriteX_62) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_7887 = _T_7885 & _T_7886; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_7888 = $signed(_T_7846) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_7889 = $signed(_T_7846) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_7890 = _T_7888 & _T_7889; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_7913 = _T_7884 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1940 = {{7'd0}, _T_7872}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_7915 = _T_7913 + _GEN_1940; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_63; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_1943 = {{1{spriteYPositionReg_63[9]}},spriteYPositionReg_63}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_7941; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_63 = _T_7941[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_7965 = {{1{inSpriteY_63[10]}},inSpriteY_63}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_7983 = inSpriteX_63; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_7991 = {{2'd0}, _T_7983}; // @[Mux.scala 80:57]
  wire [11:0] _T_7995 = {{1{inSpriteY_63[10]}},inSpriteY_63}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8003 = {{2'd0}, _T_7995}; // @[Mux.scala 80:57]
  wire  _T_8004 = $signed(inSpriteX_63) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8005 = $signed(inSpriteX_63) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8006 = _T_8004 & _T_8005; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8007 = $signed(_T_7965) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8008 = $signed(_T_7965) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8009 = _T_8007 & _T_8008; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8032 = _T_8003 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1949 = {{7'd0}, _T_7991}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8034 = _T_8032 + _GEN_1949; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_64; // @[GraphicEngineVGA.scala 355:30]
  reg [11:0] _T_8060; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_64 = _T_8060[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8084 = {{1{inSpriteY_64[10]}},inSpriteY_64}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8102 = inSpriteX_64; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8110 = {{2'd0}, _T_8102}; // @[Mux.scala 80:57]
  wire [11:0] _T_8114 = {{1{inSpriteY_64[10]}},inSpriteY_64}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8122 = {{2'd0}, _T_8114}; // @[Mux.scala 80:57]
  wire  _T_8123 = $signed(inSpriteX_64) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8124 = $signed(inSpriteX_64) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8125 = _T_8123 & _T_8124; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8126 = $signed(_T_8084) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8127 = $signed(_T_8084) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8128 = _T_8126 & _T_8127; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8151 = _T_8122 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1957 = {{7'd0}, _T_8110}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8153 = _T_8151 + _GEN_1957; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_65; // @[GraphicEngineVGA.scala 355:30]
  reg [11:0] _T_8179; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_65 = _T_8179[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8203 = {{1{inSpriteY_65[10]}},inSpriteY_65}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8221 = inSpriteX_65; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8229 = {{2'd0}, _T_8221}; // @[Mux.scala 80:57]
  wire [11:0] _T_8233 = {{1{inSpriteY_65[10]}},inSpriteY_65}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8241 = {{2'd0}, _T_8233}; // @[Mux.scala 80:57]
  wire  _T_8242 = $signed(inSpriteX_65) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8243 = $signed(inSpriteX_65) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8244 = _T_8242 & _T_8243; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8245 = $signed(_T_8203) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8246 = $signed(_T_8203) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8247 = _T_8245 & _T_8246; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8270 = _T_8241 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1965 = {{7'd0}, _T_8229}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8272 = _T_8270 + _GEN_1965; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_66; // @[GraphicEngineVGA.scala 355:30]
  reg [11:0] _T_8298; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_66 = _T_8298[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8322 = {{1{inSpriteY_66[10]}},inSpriteY_66}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8340 = inSpriteX_66; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8348 = {{2'd0}, _T_8340}; // @[Mux.scala 80:57]
  wire [11:0] _T_8352 = {{1{inSpriteY_66[10]}},inSpriteY_66}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8360 = {{2'd0}, _T_8352}; // @[Mux.scala 80:57]
  wire  _T_8361 = $signed(inSpriteX_66) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8362 = $signed(inSpriteX_66) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8363 = _T_8361 & _T_8362; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8364 = $signed(_T_8322) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8365 = $signed(_T_8322) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8366 = _T_8364 & _T_8365; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8389 = _T_8360 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1973 = {{7'd0}, _T_8348}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8391 = _T_8389 + _GEN_1973; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_67; // @[GraphicEngineVGA.scala 355:30]
  reg [11:0] _T_8417; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_67 = _T_8417[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8441 = {{1{inSpriteY_67[10]}},inSpriteY_67}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8459 = inSpriteX_67; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8467 = {{2'd0}, _T_8459}; // @[Mux.scala 80:57]
  wire [11:0] _T_8471 = {{1{inSpriteY_67[10]}},inSpriteY_67}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8479 = {{2'd0}, _T_8471}; // @[Mux.scala 80:57]
  wire  _T_8480 = $signed(inSpriteX_67) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8481 = $signed(inSpriteX_67) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8482 = _T_8480 & _T_8481; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8483 = $signed(_T_8441) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8484 = $signed(_T_8441) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8485 = _T_8483 & _T_8484; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8508 = _T_8479 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1981 = {{7'd0}, _T_8467}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8510 = _T_8508 + _GEN_1981; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_68; // @[GraphicEngineVGA.scala 355:30]
  reg [11:0] _T_8536; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_68 = _T_8536[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8560 = {{1{inSpriteY_68[10]}},inSpriteY_68}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8578 = inSpriteX_68; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8586 = {{2'd0}, _T_8578}; // @[Mux.scala 80:57]
  wire [11:0] _T_8590 = {{1{inSpriteY_68[10]}},inSpriteY_68}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8598 = {{2'd0}, _T_8590}; // @[Mux.scala 80:57]
  wire  _T_8599 = $signed(inSpriteX_68) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8600 = $signed(inSpriteX_68) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8601 = _T_8599 & _T_8600; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8602 = $signed(_T_8560) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8603 = $signed(_T_8560) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8604 = _T_8602 & _T_8603; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8627 = _T_8598 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1989 = {{7'd0}, _T_8586}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8629 = _T_8627 + _GEN_1989; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_69; // @[GraphicEngineVGA.scala 355:30]
  reg [11:0] _T_8655; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_69 = _T_8655[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8679 = {{1{inSpriteY_69[10]}},inSpriteY_69}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8697 = inSpriteX_69; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8705 = {{2'd0}, _T_8697}; // @[Mux.scala 80:57]
  wire [11:0] _T_8709 = {{1{inSpriteY_69[10]}},inSpriteY_69}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8717 = {{2'd0}, _T_8709}; // @[Mux.scala 80:57]
  wire  _T_8718 = $signed(inSpriteX_69) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8719 = $signed(inSpriteX_69) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8720 = _T_8718 & _T_8719; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8721 = $signed(_T_8679) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8722 = $signed(_T_8679) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8723 = _T_8721 & _T_8722; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8746 = _T_8717 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_1997 = {{7'd0}, _T_8705}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8748 = _T_8746 + _GEN_1997; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_70; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2000 = {{1{spriteYPositionReg_70[9]}},spriteYPositionReg_70}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_8774; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_70 = _T_8774[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8798 = {{1{inSpriteY_70[10]}},inSpriteY_70}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8816 = inSpriteX_70; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8824 = {{2'd0}, _T_8816}; // @[Mux.scala 80:57]
  wire [11:0] _T_8828 = {{1{inSpriteY_70[10]}},inSpriteY_70}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8836 = {{2'd0}, _T_8828}; // @[Mux.scala 80:57]
  wire  _T_8837 = $signed(inSpriteX_70) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8838 = $signed(inSpriteX_70) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8839 = _T_8837 & _T_8838; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8840 = $signed(_T_8798) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8841 = $signed(_T_8798) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8842 = _T_8840 & _T_8841; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8865 = _T_8836 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2006 = {{7'd0}, _T_8824}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8867 = _T_8865 + _GEN_2006; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_71; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2009 = {{1{spriteYPositionReg_71[9]}},spriteYPositionReg_71}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_8893; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_71 = _T_8893[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_8917 = {{1{inSpriteY_71[10]}},inSpriteY_71}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_8935 = inSpriteX_71; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_8943 = {{2'd0}, _T_8935}; // @[Mux.scala 80:57]
  wire [11:0] _T_8947 = {{1{inSpriteY_71[10]}},inSpriteY_71}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_8955 = {{2'd0}, _T_8947}; // @[Mux.scala 80:57]
  wire  _T_8956 = $signed(inSpriteX_71) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_8957 = $signed(inSpriteX_71) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_8958 = _T_8956 & _T_8957; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_8959 = $signed(_T_8917) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_8960 = $signed(_T_8917) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_8961 = _T_8959 & _T_8960; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_8984 = _T_8955 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2015 = {{7'd0}, _T_8943}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_8986 = _T_8984 + _GEN_2015; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_72; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2018 = {{1{spriteYPositionReg_72[9]}},spriteYPositionReg_72}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9012; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_72 = _T_9012[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9036 = {{1{inSpriteY_72[10]}},inSpriteY_72}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9054 = inSpriteX_72; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9062 = {{2'd0}, _T_9054}; // @[Mux.scala 80:57]
  wire [11:0] _T_9066 = {{1{inSpriteY_72[10]}},inSpriteY_72}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9074 = {{2'd0}, _T_9066}; // @[Mux.scala 80:57]
  wire  _T_9075 = $signed(inSpriteX_72) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9076 = $signed(inSpriteX_72) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9077 = _T_9075 & _T_9076; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9078 = $signed(_T_9036) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9079 = $signed(_T_9036) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9080 = _T_9078 & _T_9079; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9103 = _T_9074 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2024 = {{7'd0}, _T_9062}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9105 = _T_9103 + _GEN_2024; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_73; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2027 = {{1{spriteYPositionReg_73[9]}},spriteYPositionReg_73}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9131; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_73 = _T_9131[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9155 = {{1{inSpriteY_73[10]}},inSpriteY_73}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9173 = inSpriteX_73; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9181 = {{2'd0}, _T_9173}; // @[Mux.scala 80:57]
  wire [11:0] _T_9185 = {{1{inSpriteY_73[10]}},inSpriteY_73}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9193 = {{2'd0}, _T_9185}; // @[Mux.scala 80:57]
  wire  _T_9194 = $signed(inSpriteX_73) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9195 = $signed(inSpriteX_73) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9196 = _T_9194 & _T_9195; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9197 = $signed(_T_9155) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9198 = $signed(_T_9155) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9199 = _T_9197 & _T_9198; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9222 = _T_9193 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2033 = {{7'd0}, _T_9181}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9224 = _T_9222 + _GEN_2033; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_74; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2036 = {{1{spriteYPositionReg_74[9]}},spriteYPositionReg_74}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9250; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_74 = _T_9250[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9274 = {{1{inSpriteY_74[10]}},inSpriteY_74}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9292 = inSpriteX_74; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9300 = {{2'd0}, _T_9292}; // @[Mux.scala 80:57]
  wire [11:0] _T_9304 = {{1{inSpriteY_74[10]}},inSpriteY_74}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9312 = {{2'd0}, _T_9304}; // @[Mux.scala 80:57]
  wire  _T_9313 = $signed(inSpriteX_74) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9314 = $signed(inSpriteX_74) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9315 = _T_9313 & _T_9314; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9316 = $signed(_T_9274) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9317 = $signed(_T_9274) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9318 = _T_9316 & _T_9317; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9341 = _T_9312 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2042 = {{7'd0}, _T_9300}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9343 = _T_9341 + _GEN_2042; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_75; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2045 = {{1{spriteYPositionReg_75[9]}},spriteYPositionReg_75}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9369; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_75 = _T_9369[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9393 = {{1{inSpriteY_75[10]}},inSpriteY_75}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9411 = inSpriteX_75; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9419 = {{2'd0}, _T_9411}; // @[Mux.scala 80:57]
  wire [11:0] _T_9423 = {{1{inSpriteY_75[10]}},inSpriteY_75}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9431 = {{2'd0}, _T_9423}; // @[Mux.scala 80:57]
  wire  _T_9432 = $signed(inSpriteX_75) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9433 = $signed(inSpriteX_75) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9434 = _T_9432 & _T_9433; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9435 = $signed(_T_9393) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9436 = $signed(_T_9393) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9437 = _T_9435 & _T_9436; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9460 = _T_9431 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2051 = {{7'd0}, _T_9419}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9462 = _T_9460 + _GEN_2051; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_76; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2054 = {{1{spriteYPositionReg_76[9]}},spriteYPositionReg_76}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9488; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_76 = _T_9488[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9512 = {{1{inSpriteY_76[10]}},inSpriteY_76}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9530 = inSpriteX_76; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9538 = {{2'd0}, _T_9530}; // @[Mux.scala 80:57]
  wire [11:0] _T_9542 = {{1{inSpriteY_76[10]}},inSpriteY_76}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9550 = {{2'd0}, _T_9542}; // @[Mux.scala 80:57]
  wire  _T_9551 = $signed(inSpriteX_76) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9552 = $signed(inSpriteX_76) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9553 = _T_9551 & _T_9552; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9554 = $signed(_T_9512) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9555 = $signed(_T_9512) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9556 = _T_9554 & _T_9555; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9579 = _T_9550 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2060 = {{7'd0}, _T_9538}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9581 = _T_9579 + _GEN_2060; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_77; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2063 = {{1{spriteYPositionReg_77[9]}},spriteYPositionReg_77}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9607; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_77 = _T_9607[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9631 = {{1{inSpriteY_77[10]}},inSpriteY_77}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9649 = inSpriteX_77; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9657 = {{2'd0}, _T_9649}; // @[Mux.scala 80:57]
  wire [11:0] _T_9661 = {{1{inSpriteY_77[10]}},inSpriteY_77}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9669 = {{2'd0}, _T_9661}; // @[Mux.scala 80:57]
  wire  _T_9670 = $signed(inSpriteX_77) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9671 = $signed(inSpriteX_77) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9672 = _T_9670 & _T_9671; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9673 = $signed(_T_9631) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9674 = $signed(_T_9631) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9675 = _T_9673 & _T_9674; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9698 = _T_9669 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2069 = {{7'd0}, _T_9657}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9700 = _T_9698 + _GEN_2069; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_78; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2072 = {{1{spriteYPositionReg_78[9]}},spriteYPositionReg_78}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9726; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_78 = _T_9726[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9750 = {{1{inSpriteY_78[10]}},inSpriteY_78}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9768 = inSpriteX_78; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9776 = {{2'd0}, _T_9768}; // @[Mux.scala 80:57]
  wire [11:0] _T_9780 = {{1{inSpriteY_78[10]}},inSpriteY_78}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9788 = {{2'd0}, _T_9780}; // @[Mux.scala 80:57]
  wire  _T_9789 = $signed(inSpriteX_78) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9790 = $signed(inSpriteX_78) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9791 = _T_9789 & _T_9790; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9792 = $signed(_T_9750) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9793 = $signed(_T_9750) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9794 = _T_9792 & _T_9793; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9817 = _T_9788 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2078 = {{7'd0}, _T_9776}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9819 = _T_9817 + _GEN_2078; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_79; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2081 = {{1{spriteYPositionReg_79[9]}},spriteYPositionReg_79}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9845; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_79 = _T_9845[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9869 = {{1{inSpriteY_79[10]}},inSpriteY_79}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_9887 = inSpriteX_79; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_9895 = {{2'd0}, _T_9887}; // @[Mux.scala 80:57]
  wire [11:0] _T_9899 = {{1{inSpriteY_79[10]}},inSpriteY_79}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_9907 = {{2'd0}, _T_9899}; // @[Mux.scala 80:57]
  wire  _T_9908 = $signed(inSpriteX_79) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_9909 = $signed(inSpriteX_79) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_9910 = _T_9908 & _T_9909; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_9911 = $signed(_T_9869) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_9912 = $signed(_T_9869) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_9913 = _T_9911 & _T_9912; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_9936 = _T_9907 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2087 = {{7'd0}, _T_9895}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_9938 = _T_9936 + _GEN_2087; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_80; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2090 = {{1{spriteYPositionReg_80[9]}},spriteYPositionReg_80}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_9964; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_80 = _T_9964[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_9988 = {{1{inSpriteY_80[10]}},inSpriteY_80}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10006 = inSpriteX_80; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10014 = {{2'd0}, _T_10006}; // @[Mux.scala 80:57]
  wire [11:0] _T_10018 = {{1{inSpriteY_80[10]}},inSpriteY_80}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10026 = {{2'd0}, _T_10018}; // @[Mux.scala 80:57]
  wire  _T_10027 = $signed(inSpriteX_80) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10028 = $signed(inSpriteX_80) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10029 = _T_10027 & _T_10028; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10030 = $signed(_T_9988) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10031 = $signed(_T_9988) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10032 = _T_10030 & _T_10031; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10055 = _T_10026 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2096 = {{7'd0}, _T_10014}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10057 = _T_10055 + _GEN_2096; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_81; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2099 = {{1{spriteYPositionReg_81[9]}},spriteYPositionReg_81}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10083; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_81 = _T_10083[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10107 = {{1{inSpriteY_81[10]}},inSpriteY_81}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10125 = inSpriteX_81; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10133 = {{2'd0}, _T_10125}; // @[Mux.scala 80:57]
  wire [11:0] _T_10137 = {{1{inSpriteY_81[10]}},inSpriteY_81}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10145 = {{2'd0}, _T_10137}; // @[Mux.scala 80:57]
  wire  _T_10146 = $signed(inSpriteX_81) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10147 = $signed(inSpriteX_81) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10148 = _T_10146 & _T_10147; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10149 = $signed(_T_10107) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10150 = $signed(_T_10107) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10151 = _T_10149 & _T_10150; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10174 = _T_10145 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2105 = {{7'd0}, _T_10133}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10176 = _T_10174 + _GEN_2105; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_82; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2108 = {{1{spriteYPositionReg_82[9]}},spriteYPositionReg_82}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10202; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_82 = _T_10202[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10226 = {{1{inSpriteY_82[10]}},inSpriteY_82}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10244 = inSpriteX_82; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10252 = {{2'd0}, _T_10244}; // @[Mux.scala 80:57]
  wire [11:0] _T_10256 = {{1{inSpriteY_82[10]}},inSpriteY_82}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10264 = {{2'd0}, _T_10256}; // @[Mux.scala 80:57]
  wire  _T_10265 = $signed(inSpriteX_82) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10266 = $signed(inSpriteX_82) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10267 = _T_10265 & _T_10266; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10268 = $signed(_T_10226) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10269 = $signed(_T_10226) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10270 = _T_10268 & _T_10269; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10293 = _T_10264 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2114 = {{7'd0}, _T_10252}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10295 = _T_10293 + _GEN_2114; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_83; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2117 = {{1{spriteYPositionReg_83[9]}},spriteYPositionReg_83}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10321; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_83 = _T_10321[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10345 = {{1{inSpriteY_83[10]}},inSpriteY_83}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10363 = inSpriteX_83; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10371 = {{2'd0}, _T_10363}; // @[Mux.scala 80:57]
  wire [11:0] _T_10375 = {{1{inSpriteY_83[10]}},inSpriteY_83}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10383 = {{2'd0}, _T_10375}; // @[Mux.scala 80:57]
  wire  _T_10384 = $signed(inSpriteX_83) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10385 = $signed(inSpriteX_83) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10386 = _T_10384 & _T_10385; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10387 = $signed(_T_10345) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10388 = $signed(_T_10345) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10389 = _T_10387 & _T_10388; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10412 = _T_10383 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2123 = {{7'd0}, _T_10371}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10414 = _T_10412 + _GEN_2123; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_84; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2126 = {{1{spriteYPositionReg_84[9]}},spriteYPositionReg_84}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10440; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_84 = _T_10440[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10464 = {{1{inSpriteY_84[10]}},inSpriteY_84}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10482 = inSpriteX_84; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10490 = {{2'd0}, _T_10482}; // @[Mux.scala 80:57]
  wire [11:0] _T_10494 = {{1{inSpriteY_84[10]}},inSpriteY_84}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10502 = {{2'd0}, _T_10494}; // @[Mux.scala 80:57]
  wire  _T_10503 = $signed(inSpriteX_84) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10504 = $signed(inSpriteX_84) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10505 = _T_10503 & _T_10504; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10506 = $signed(_T_10464) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10507 = $signed(_T_10464) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10508 = _T_10506 & _T_10507; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10531 = _T_10502 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2132 = {{7'd0}, _T_10490}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10533 = _T_10531 + _GEN_2132; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_85; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2135 = {{1{spriteYPositionReg_85[9]}},spriteYPositionReg_85}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10559; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_85 = _T_10559[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10583 = {{1{inSpriteY_85[10]}},inSpriteY_85}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10601 = inSpriteX_85; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10609 = {{2'd0}, _T_10601}; // @[Mux.scala 80:57]
  wire [11:0] _T_10613 = {{1{inSpriteY_85[10]}},inSpriteY_85}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10621 = {{2'd0}, _T_10613}; // @[Mux.scala 80:57]
  wire  _T_10622 = $signed(inSpriteX_85) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10623 = $signed(inSpriteX_85) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10624 = _T_10622 & _T_10623; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10625 = $signed(_T_10583) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10626 = $signed(_T_10583) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10627 = _T_10625 & _T_10626; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10650 = _T_10621 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2141 = {{7'd0}, _T_10609}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10652 = _T_10650 + _GEN_2141; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_86; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2144 = {{1{spriteYPositionReg_86[9]}},spriteYPositionReg_86}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10678; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_86 = _T_10678[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10702 = {{1{inSpriteY_86[10]}},inSpriteY_86}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10720 = inSpriteX_86; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10728 = {{2'd0}, _T_10720}; // @[Mux.scala 80:57]
  wire [11:0] _T_10732 = {{1{inSpriteY_86[10]}},inSpriteY_86}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10740 = {{2'd0}, _T_10732}; // @[Mux.scala 80:57]
  wire  _T_10741 = $signed(inSpriteX_86) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10742 = $signed(inSpriteX_86) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10743 = _T_10741 & _T_10742; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10744 = $signed(_T_10702) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10745 = $signed(_T_10702) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10746 = _T_10744 & _T_10745; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10769 = _T_10740 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2150 = {{7'd0}, _T_10728}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10771 = _T_10769 + _GEN_2150; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_87; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2153 = {{1{spriteYPositionReg_87[9]}},spriteYPositionReg_87}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10797; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_87 = _T_10797[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10821 = {{1{inSpriteY_87[10]}},inSpriteY_87}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10839 = inSpriteX_87; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10847 = {{2'd0}, _T_10839}; // @[Mux.scala 80:57]
  wire [11:0] _T_10851 = {{1{inSpriteY_87[10]}},inSpriteY_87}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10859 = {{2'd0}, _T_10851}; // @[Mux.scala 80:57]
  wire  _T_10860 = $signed(inSpriteX_87) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10861 = $signed(inSpriteX_87) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10862 = _T_10860 & _T_10861; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10863 = $signed(_T_10821) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10864 = $signed(_T_10821) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10865 = _T_10863 & _T_10864; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_10888 = _T_10859 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2159 = {{7'd0}, _T_10847}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_10890 = _T_10888 + _GEN_2159; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_88; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2162 = {{1{spriteYPositionReg_88[9]}},spriteYPositionReg_88}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_10916; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_88 = _T_10916[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_10940 = {{1{inSpriteY_88[10]}},inSpriteY_88}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_10958 = inSpriteX_88; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_10966 = {{2'd0}, _T_10958}; // @[Mux.scala 80:57]
  wire [11:0] _T_10970 = {{1{inSpriteY_88[10]}},inSpriteY_88}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_10978 = {{2'd0}, _T_10970}; // @[Mux.scala 80:57]
  wire  _T_10979 = $signed(inSpriteX_88) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_10980 = $signed(inSpriteX_88) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_10981 = _T_10979 & _T_10980; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_10982 = $signed(_T_10940) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_10983 = $signed(_T_10940) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_10984 = _T_10982 & _T_10983; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11007 = _T_10978 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2168 = {{7'd0}, _T_10966}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11009 = _T_11007 + _GEN_2168; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_89; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2171 = {{1{spriteYPositionReg_89[9]}},spriteYPositionReg_89}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11035; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_89 = _T_11035[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11059 = {{1{inSpriteY_89[10]}},inSpriteY_89}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11077 = inSpriteX_89; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11085 = {{2'd0}, _T_11077}; // @[Mux.scala 80:57]
  wire [11:0] _T_11089 = {{1{inSpriteY_89[10]}},inSpriteY_89}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11097 = {{2'd0}, _T_11089}; // @[Mux.scala 80:57]
  wire  _T_11098 = $signed(inSpriteX_89) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11099 = $signed(inSpriteX_89) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11100 = _T_11098 & _T_11099; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11101 = $signed(_T_11059) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11102 = $signed(_T_11059) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11103 = _T_11101 & _T_11102; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11126 = _T_11097 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2177 = {{7'd0}, _T_11085}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11128 = _T_11126 + _GEN_2177; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_90; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2180 = {{1{spriteYPositionReg_90[9]}},spriteYPositionReg_90}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11154; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_90 = _T_11154[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11178 = {{1{inSpriteY_90[10]}},inSpriteY_90}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11196 = inSpriteX_90; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11204 = {{2'd0}, _T_11196}; // @[Mux.scala 80:57]
  wire [11:0] _T_11208 = {{1{inSpriteY_90[10]}},inSpriteY_90}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11216 = {{2'd0}, _T_11208}; // @[Mux.scala 80:57]
  wire  _T_11217 = $signed(inSpriteX_90) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11218 = $signed(inSpriteX_90) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11219 = _T_11217 & _T_11218; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11220 = $signed(_T_11178) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11221 = $signed(_T_11178) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11222 = _T_11220 & _T_11221; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11245 = _T_11216 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2186 = {{7'd0}, _T_11204}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11247 = _T_11245 + _GEN_2186; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_91; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2189 = {{1{spriteYPositionReg_91[9]}},spriteYPositionReg_91}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11273; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_91 = _T_11273[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11297 = {{1{inSpriteY_91[10]}},inSpriteY_91}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11315 = inSpriteX_91; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11323 = {{2'd0}, _T_11315}; // @[Mux.scala 80:57]
  wire [11:0] _T_11327 = {{1{inSpriteY_91[10]}},inSpriteY_91}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11335 = {{2'd0}, _T_11327}; // @[Mux.scala 80:57]
  wire  _T_11336 = $signed(inSpriteX_91) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11337 = $signed(inSpriteX_91) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11338 = _T_11336 & _T_11337; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11339 = $signed(_T_11297) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11340 = $signed(_T_11297) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11341 = _T_11339 & _T_11340; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11364 = _T_11335 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2195 = {{7'd0}, _T_11323}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11366 = _T_11364 + _GEN_2195; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_92; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2198 = {{1{spriteYPositionReg_92[9]}},spriteYPositionReg_92}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11392; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_92 = _T_11392[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11416 = {{1{inSpriteY_92[10]}},inSpriteY_92}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11434 = inSpriteX_92; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11442 = {{2'd0}, _T_11434}; // @[Mux.scala 80:57]
  wire [11:0] _T_11446 = {{1{inSpriteY_92[10]}},inSpriteY_92}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11454 = {{2'd0}, _T_11446}; // @[Mux.scala 80:57]
  wire  _T_11455 = $signed(inSpriteX_92) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11456 = $signed(inSpriteX_92) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11457 = _T_11455 & _T_11456; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11458 = $signed(_T_11416) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11459 = $signed(_T_11416) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11460 = _T_11458 & _T_11459; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11483 = _T_11454 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2204 = {{7'd0}, _T_11442}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11485 = _T_11483 + _GEN_2204; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_93; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2207 = {{1{spriteYPositionReg_93[9]}},spriteYPositionReg_93}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11511; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_93 = _T_11511[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11535 = {{1{inSpriteY_93[10]}},inSpriteY_93}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11553 = inSpriteX_93; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11561 = {{2'd0}, _T_11553}; // @[Mux.scala 80:57]
  wire [11:0] _T_11565 = {{1{inSpriteY_93[10]}},inSpriteY_93}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11573 = {{2'd0}, _T_11565}; // @[Mux.scala 80:57]
  wire  _T_11574 = $signed(inSpriteX_93) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11575 = $signed(inSpriteX_93) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11576 = _T_11574 & _T_11575; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11577 = $signed(_T_11535) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11578 = $signed(_T_11535) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11579 = _T_11577 & _T_11578; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11602 = _T_11573 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2213 = {{7'd0}, _T_11561}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11604 = _T_11602 + _GEN_2213; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_94; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2216 = {{1{spriteYPositionReg_94[9]}},spriteYPositionReg_94}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11630; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_94 = _T_11630[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11654 = {{1{inSpriteY_94[10]}},inSpriteY_94}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11672 = inSpriteX_94; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11680 = {{2'd0}, _T_11672}; // @[Mux.scala 80:57]
  wire [11:0] _T_11684 = {{1{inSpriteY_94[10]}},inSpriteY_94}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11692 = {{2'd0}, _T_11684}; // @[Mux.scala 80:57]
  wire  _T_11693 = $signed(inSpriteX_94) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11694 = $signed(inSpriteX_94) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11695 = _T_11693 & _T_11694; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11696 = $signed(_T_11654) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11697 = $signed(_T_11654) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11698 = _T_11696 & _T_11697; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11721 = _T_11692 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2222 = {{7'd0}, _T_11680}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11723 = _T_11721 + _GEN_2222; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_95; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2225 = {{1{spriteYPositionReg_95[9]}},spriteYPositionReg_95}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11749; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_95 = _T_11749[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11773 = {{1{inSpriteY_95[10]}},inSpriteY_95}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11791 = inSpriteX_95; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11799 = {{2'd0}, _T_11791}; // @[Mux.scala 80:57]
  wire [11:0] _T_11803 = {{1{inSpriteY_95[10]}},inSpriteY_95}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11811 = {{2'd0}, _T_11803}; // @[Mux.scala 80:57]
  wire  _T_11812 = $signed(inSpriteX_95) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11813 = $signed(inSpriteX_95) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11814 = _T_11812 & _T_11813; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11815 = $signed(_T_11773) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11816 = $signed(_T_11773) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11817 = _T_11815 & _T_11816; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11840 = _T_11811 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2231 = {{7'd0}, _T_11799}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11842 = _T_11840 + _GEN_2231; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_96; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2234 = {{1{spriteYPositionReg_96[9]}},spriteYPositionReg_96}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11868; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_96 = _T_11868[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_11892 = {{1{inSpriteY_96[10]}},inSpriteY_96}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_11910 = inSpriteX_96; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_11918 = {{2'd0}, _T_11910}; // @[Mux.scala 80:57]
  wire [11:0] _T_11922 = {{1{inSpriteY_96[10]}},inSpriteY_96}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_11930 = {{2'd0}, _T_11922}; // @[Mux.scala 80:57]
  wire  _T_11931 = $signed(inSpriteX_96) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_11932 = $signed(inSpriteX_96) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_11933 = _T_11931 & _T_11932; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_11934 = $signed(_T_11892) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_11935 = $signed(_T_11892) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_11936 = _T_11934 & _T_11935; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_11959 = _T_11930 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2240 = {{7'd0}, _T_11918}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_11961 = _T_11959 + _GEN_2240; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_97; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2243 = {{1{spriteYPositionReg_97[9]}},spriteYPositionReg_97}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_11987; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_97 = _T_11987[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12011 = {{1{inSpriteY_97[10]}},inSpriteY_97}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12029 = inSpriteX_97; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12037 = {{2'd0}, _T_12029}; // @[Mux.scala 80:57]
  wire [11:0] _T_12041 = {{1{inSpriteY_97[10]}},inSpriteY_97}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12049 = {{2'd0}, _T_12041}; // @[Mux.scala 80:57]
  wire  _T_12050 = $signed(inSpriteX_97) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12051 = $signed(inSpriteX_97) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12052 = _T_12050 & _T_12051; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12053 = $signed(_T_12011) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12054 = $signed(_T_12011) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12055 = _T_12053 & _T_12054; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12078 = _T_12049 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2249 = {{7'd0}, _T_12037}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12080 = _T_12078 + _GEN_2249; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_98; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2252 = {{1{spriteYPositionReg_98[9]}},spriteYPositionReg_98}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12106; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_98 = _T_12106[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12130 = {{1{inSpriteY_98[10]}},inSpriteY_98}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12148 = inSpriteX_98; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12156 = {{2'd0}, _T_12148}; // @[Mux.scala 80:57]
  wire [11:0] _T_12160 = {{1{inSpriteY_98[10]}},inSpriteY_98}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12168 = {{2'd0}, _T_12160}; // @[Mux.scala 80:57]
  wire  _T_12169 = $signed(inSpriteX_98) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12170 = $signed(inSpriteX_98) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12171 = _T_12169 & _T_12170; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12172 = $signed(_T_12130) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12173 = $signed(_T_12130) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12174 = _T_12172 & _T_12173; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12197 = _T_12168 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2258 = {{7'd0}, _T_12156}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12199 = _T_12197 + _GEN_2258; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_99; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2261 = {{1{spriteYPositionReg_99[9]}},spriteYPositionReg_99}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12225; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_99 = _T_12225[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12249 = {{1{inSpriteY_99[10]}},inSpriteY_99}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12267 = inSpriteX_99; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12275 = {{2'd0}, _T_12267}; // @[Mux.scala 80:57]
  wire [11:0] _T_12279 = {{1{inSpriteY_99[10]}},inSpriteY_99}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12287 = {{2'd0}, _T_12279}; // @[Mux.scala 80:57]
  wire  _T_12288 = $signed(inSpriteX_99) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12289 = $signed(inSpriteX_99) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12290 = _T_12288 & _T_12289; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12291 = $signed(_T_12249) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12292 = $signed(_T_12249) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12293 = _T_12291 & _T_12292; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12316 = _T_12287 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2267 = {{7'd0}, _T_12275}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12318 = _T_12316 + _GEN_2267; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_100; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2270 = {{1{spriteYPositionReg_100[9]}},spriteYPositionReg_100}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12344; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_100 = _T_12344[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12368 = {{1{inSpriteY_100[10]}},inSpriteY_100}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12386 = inSpriteX_100; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12394 = {{2'd0}, _T_12386}; // @[Mux.scala 80:57]
  wire [11:0] _T_12398 = {{1{inSpriteY_100[10]}},inSpriteY_100}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12406 = {{2'd0}, _T_12398}; // @[Mux.scala 80:57]
  wire  _T_12407 = $signed(inSpriteX_100) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12408 = $signed(inSpriteX_100) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12409 = _T_12407 & _T_12408; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12410 = $signed(_T_12368) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12411 = $signed(_T_12368) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12412 = _T_12410 & _T_12411; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12435 = _T_12406 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2276 = {{7'd0}, _T_12394}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12437 = _T_12435 + _GEN_2276; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_101; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2279 = {{1{spriteYPositionReg_101[9]}},spriteYPositionReg_101}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12463; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_101 = _T_12463[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12487 = {{1{inSpriteY_101[10]}},inSpriteY_101}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12505 = inSpriteX_101; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12513 = {{2'd0}, _T_12505}; // @[Mux.scala 80:57]
  wire [11:0] _T_12517 = {{1{inSpriteY_101[10]}},inSpriteY_101}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12525 = {{2'd0}, _T_12517}; // @[Mux.scala 80:57]
  wire  _T_12526 = $signed(inSpriteX_101) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12527 = $signed(inSpriteX_101) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12528 = _T_12526 & _T_12527; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12529 = $signed(_T_12487) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12530 = $signed(_T_12487) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12531 = _T_12529 & _T_12530; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12554 = _T_12525 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2285 = {{7'd0}, _T_12513}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12556 = _T_12554 + _GEN_2285; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_102; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2288 = {{1{spriteYPositionReg_102[9]}},spriteYPositionReg_102}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12582; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_102 = _T_12582[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12606 = {{1{inSpriteY_102[10]}},inSpriteY_102}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12624 = inSpriteX_102; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12632 = {{2'd0}, _T_12624}; // @[Mux.scala 80:57]
  wire [11:0] _T_12636 = {{1{inSpriteY_102[10]}},inSpriteY_102}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12644 = {{2'd0}, _T_12636}; // @[Mux.scala 80:57]
  wire  _T_12645 = $signed(inSpriteX_102) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12646 = $signed(inSpriteX_102) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12647 = _T_12645 & _T_12646; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12648 = $signed(_T_12606) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12649 = $signed(_T_12606) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12650 = _T_12648 & _T_12649; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12673 = _T_12644 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2294 = {{7'd0}, _T_12632}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12675 = _T_12673 + _GEN_2294; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_103; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2297 = {{1{spriteYPositionReg_103[9]}},spriteYPositionReg_103}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12701; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_103 = _T_12701[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12725 = {{1{inSpriteY_103[10]}},inSpriteY_103}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12743 = inSpriteX_103; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12751 = {{2'd0}, _T_12743}; // @[Mux.scala 80:57]
  wire [11:0] _T_12755 = {{1{inSpriteY_103[10]}},inSpriteY_103}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12763 = {{2'd0}, _T_12755}; // @[Mux.scala 80:57]
  wire  _T_12764 = $signed(inSpriteX_103) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12765 = $signed(inSpriteX_103) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12766 = _T_12764 & _T_12765; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12767 = $signed(_T_12725) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12768 = $signed(_T_12725) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12769 = _T_12767 & _T_12768; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12792 = _T_12763 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2303 = {{7'd0}, _T_12751}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12794 = _T_12792 + _GEN_2303; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_104; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2306 = {{1{spriteYPositionReg_104[9]}},spriteYPositionReg_104}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12820; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_104 = _T_12820[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12844 = {{1{inSpriteY_104[10]}},inSpriteY_104}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12862 = inSpriteX_104; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12870 = {{2'd0}, _T_12862}; // @[Mux.scala 80:57]
  wire [11:0] _T_12874 = {{1{inSpriteY_104[10]}},inSpriteY_104}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_12882 = {{2'd0}, _T_12874}; // @[Mux.scala 80:57]
  wire  _T_12883 = $signed(inSpriteX_104) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_12884 = $signed(inSpriteX_104) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_12885 = _T_12883 & _T_12884; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_12886 = $signed(_T_12844) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_12887 = $signed(_T_12844) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_12888 = _T_12886 & _T_12887; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_12911 = _T_12882 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2312 = {{7'd0}, _T_12870}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_12913 = _T_12911 + _GEN_2312; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_105; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2315 = {{1{spriteYPositionReg_105[9]}},spriteYPositionReg_105}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_12939; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_105 = _T_12939[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_12963 = {{1{inSpriteY_105[10]}},inSpriteY_105}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_12981 = inSpriteX_105; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_12989 = {{2'd0}, _T_12981}; // @[Mux.scala 80:57]
  wire [11:0] _T_12993 = {{1{inSpriteY_105[10]}},inSpriteY_105}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13001 = {{2'd0}, _T_12993}; // @[Mux.scala 80:57]
  wire  _T_13002 = $signed(inSpriteX_105) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13003 = $signed(inSpriteX_105) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13004 = _T_13002 & _T_13003; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13005 = $signed(_T_12963) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13006 = $signed(_T_12963) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13007 = _T_13005 & _T_13006; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13030 = _T_13001 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2321 = {{7'd0}, _T_12989}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13032 = _T_13030 + _GEN_2321; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_106; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2324 = {{1{spriteYPositionReg_106[9]}},spriteYPositionReg_106}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13058; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_106 = _T_13058[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13082 = {{1{inSpriteY_106[10]}},inSpriteY_106}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13100 = inSpriteX_106; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13108 = {{2'd0}, _T_13100}; // @[Mux.scala 80:57]
  wire [11:0] _T_13112 = {{1{inSpriteY_106[10]}},inSpriteY_106}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13120 = {{2'd0}, _T_13112}; // @[Mux.scala 80:57]
  wire  _T_13121 = $signed(inSpriteX_106) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13122 = $signed(inSpriteX_106) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13123 = _T_13121 & _T_13122; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13124 = $signed(_T_13082) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13125 = $signed(_T_13082) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13126 = _T_13124 & _T_13125; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13149 = _T_13120 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2330 = {{7'd0}, _T_13108}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13151 = _T_13149 + _GEN_2330; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_107; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2333 = {{1{spriteYPositionReg_107[9]}},spriteYPositionReg_107}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13177; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_107 = _T_13177[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13201 = {{1{inSpriteY_107[10]}},inSpriteY_107}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13219 = inSpriteX_107; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13227 = {{2'd0}, _T_13219}; // @[Mux.scala 80:57]
  wire [11:0] _T_13231 = {{1{inSpriteY_107[10]}},inSpriteY_107}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13239 = {{2'd0}, _T_13231}; // @[Mux.scala 80:57]
  wire  _T_13240 = $signed(inSpriteX_107) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13241 = $signed(inSpriteX_107) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13242 = _T_13240 & _T_13241; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13243 = $signed(_T_13201) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13244 = $signed(_T_13201) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13245 = _T_13243 & _T_13244; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13268 = _T_13239 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2339 = {{7'd0}, _T_13227}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13270 = _T_13268 + _GEN_2339; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_108; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2342 = {{1{spriteYPositionReg_108[9]}},spriteYPositionReg_108}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13296; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_108 = _T_13296[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13320 = {{1{inSpriteY_108[10]}},inSpriteY_108}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13338 = inSpriteX_108; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13346 = {{2'd0}, _T_13338}; // @[Mux.scala 80:57]
  wire [11:0] _T_13350 = {{1{inSpriteY_108[10]}},inSpriteY_108}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13358 = {{2'd0}, _T_13350}; // @[Mux.scala 80:57]
  wire  _T_13359 = $signed(inSpriteX_108) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13360 = $signed(inSpriteX_108) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13361 = _T_13359 & _T_13360; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13362 = $signed(_T_13320) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13363 = $signed(_T_13320) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13364 = _T_13362 & _T_13363; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13387 = _T_13358 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2348 = {{7'd0}, _T_13346}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13389 = _T_13387 + _GEN_2348; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_109; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2351 = {{1{spriteYPositionReg_109[9]}},spriteYPositionReg_109}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13415; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_109 = _T_13415[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13439 = {{1{inSpriteY_109[10]}},inSpriteY_109}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13457 = inSpriteX_109; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13465 = {{2'd0}, _T_13457}; // @[Mux.scala 80:57]
  wire [11:0] _T_13469 = {{1{inSpriteY_109[10]}},inSpriteY_109}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13477 = {{2'd0}, _T_13469}; // @[Mux.scala 80:57]
  wire  _T_13478 = $signed(inSpriteX_109) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13479 = $signed(inSpriteX_109) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13480 = _T_13478 & _T_13479; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13481 = $signed(_T_13439) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13482 = $signed(_T_13439) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13483 = _T_13481 & _T_13482; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13506 = _T_13477 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2357 = {{7'd0}, _T_13465}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13508 = _T_13506 + _GEN_2357; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_110; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2360 = {{1{spriteYPositionReg_110[9]}},spriteYPositionReg_110}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13534; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_110 = _T_13534[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13558 = {{1{inSpriteY_110[10]}},inSpriteY_110}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13576 = inSpriteX_110; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13584 = {{2'd0}, _T_13576}; // @[Mux.scala 80:57]
  wire [11:0] _T_13588 = {{1{inSpriteY_110[10]}},inSpriteY_110}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13596 = {{2'd0}, _T_13588}; // @[Mux.scala 80:57]
  wire  _T_13597 = $signed(inSpriteX_110) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13598 = $signed(inSpriteX_110) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13599 = _T_13597 & _T_13598; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13600 = $signed(_T_13558) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13601 = $signed(_T_13558) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13602 = _T_13600 & _T_13601; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13625 = _T_13596 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2366 = {{7'd0}, _T_13584}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13627 = _T_13625 + _GEN_2366; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_111; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2369 = {{1{spriteYPositionReg_111[9]}},spriteYPositionReg_111}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13653; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_111 = _T_13653[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13677 = {{1{inSpriteY_111[10]}},inSpriteY_111}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13695 = inSpriteX_111; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13703 = {{2'd0}, _T_13695}; // @[Mux.scala 80:57]
  wire [11:0] _T_13707 = {{1{inSpriteY_111[10]}},inSpriteY_111}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13715 = {{2'd0}, _T_13707}; // @[Mux.scala 80:57]
  wire  _T_13716 = $signed(inSpriteX_111) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13717 = $signed(inSpriteX_111) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13718 = _T_13716 & _T_13717; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13719 = $signed(_T_13677) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13720 = $signed(_T_13677) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13721 = _T_13719 & _T_13720; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13744 = _T_13715 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2375 = {{7'd0}, _T_13703}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13746 = _T_13744 + _GEN_2375; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_112; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2378 = {{1{spriteYPositionReg_112[9]}},spriteYPositionReg_112}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13772; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_112 = _T_13772[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13796 = {{1{inSpriteY_112[10]}},inSpriteY_112}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13814 = inSpriteX_112; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13822 = {{2'd0}, _T_13814}; // @[Mux.scala 80:57]
  wire [11:0] _T_13826 = {{1{inSpriteY_112[10]}},inSpriteY_112}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13834 = {{2'd0}, _T_13826}; // @[Mux.scala 80:57]
  wire  _T_13835 = $signed(inSpriteX_112) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13836 = $signed(inSpriteX_112) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13837 = _T_13835 & _T_13836; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13838 = $signed(_T_13796) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13839 = $signed(_T_13796) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13840 = _T_13838 & _T_13839; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13863 = _T_13834 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2384 = {{7'd0}, _T_13822}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13865 = _T_13863 + _GEN_2384; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_113; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2387 = {{1{spriteYPositionReg_113[9]}},spriteYPositionReg_113}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_13891; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_113 = _T_13891[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_13915 = {{1{inSpriteY_113[10]}},inSpriteY_113}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_13933 = inSpriteX_113; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_13941 = {{2'd0}, _T_13933}; // @[Mux.scala 80:57]
  wire [11:0] _T_13945 = {{1{inSpriteY_113[10]}},inSpriteY_113}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_13953 = {{2'd0}, _T_13945}; // @[Mux.scala 80:57]
  wire  _T_13954 = $signed(inSpriteX_113) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_13955 = $signed(inSpriteX_113) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_13956 = _T_13954 & _T_13955; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_13957 = $signed(_T_13915) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_13958 = $signed(_T_13915) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_13959 = _T_13957 & _T_13958; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_13982 = _T_13953 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2393 = {{7'd0}, _T_13941}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_13984 = _T_13982 + _GEN_2393; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_114; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2396 = {{1{spriteYPositionReg_114[9]}},spriteYPositionReg_114}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14010; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_114 = _T_14010[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14034 = {{1{inSpriteY_114[10]}},inSpriteY_114}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14052 = inSpriteX_114; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14060 = {{2'd0}, _T_14052}; // @[Mux.scala 80:57]
  wire [11:0] _T_14064 = {{1{inSpriteY_114[10]}},inSpriteY_114}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14072 = {{2'd0}, _T_14064}; // @[Mux.scala 80:57]
  wire  _T_14073 = $signed(inSpriteX_114) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14074 = $signed(inSpriteX_114) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14075 = _T_14073 & _T_14074; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14076 = $signed(_T_14034) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14077 = $signed(_T_14034) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14078 = _T_14076 & _T_14077; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14101 = _T_14072 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2402 = {{7'd0}, _T_14060}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14103 = _T_14101 + _GEN_2402; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_115; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2405 = {{1{spriteYPositionReg_115[9]}},spriteYPositionReg_115}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14129; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_115 = _T_14129[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14153 = {{1{inSpriteY_115[10]}},inSpriteY_115}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14171 = inSpriteX_115; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14179 = {{2'd0}, _T_14171}; // @[Mux.scala 80:57]
  wire [11:0] _T_14183 = {{1{inSpriteY_115[10]}},inSpriteY_115}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14191 = {{2'd0}, _T_14183}; // @[Mux.scala 80:57]
  wire  _T_14192 = $signed(inSpriteX_115) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14193 = $signed(inSpriteX_115) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14194 = _T_14192 & _T_14193; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14195 = $signed(_T_14153) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14196 = $signed(_T_14153) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14197 = _T_14195 & _T_14196; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14220 = _T_14191 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2411 = {{7'd0}, _T_14179}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14222 = _T_14220 + _GEN_2411; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_116; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2414 = {{1{spriteYPositionReg_116[9]}},spriteYPositionReg_116}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14248; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_116 = _T_14248[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14272 = {{1{inSpriteY_116[10]}},inSpriteY_116}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14290 = inSpriteX_116; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14298 = {{2'd0}, _T_14290}; // @[Mux.scala 80:57]
  wire [11:0] _T_14302 = {{1{inSpriteY_116[10]}},inSpriteY_116}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14310 = {{2'd0}, _T_14302}; // @[Mux.scala 80:57]
  wire  _T_14311 = $signed(inSpriteX_116) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14312 = $signed(inSpriteX_116) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14313 = _T_14311 & _T_14312; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14314 = $signed(_T_14272) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14315 = $signed(_T_14272) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14316 = _T_14314 & _T_14315; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14339 = _T_14310 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2420 = {{7'd0}, _T_14298}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14341 = _T_14339 + _GEN_2420; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_117; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2423 = {{1{spriteYPositionReg_117[9]}},spriteYPositionReg_117}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14367; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_117 = _T_14367[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14391 = {{1{inSpriteY_117[10]}},inSpriteY_117}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14409 = inSpriteX_117; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14417 = {{2'd0}, _T_14409}; // @[Mux.scala 80:57]
  wire [11:0] _T_14421 = {{1{inSpriteY_117[10]}},inSpriteY_117}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14429 = {{2'd0}, _T_14421}; // @[Mux.scala 80:57]
  wire  _T_14430 = $signed(inSpriteX_117) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14431 = $signed(inSpriteX_117) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14432 = _T_14430 & _T_14431; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14433 = $signed(_T_14391) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14434 = $signed(_T_14391) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14435 = _T_14433 & _T_14434; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14458 = _T_14429 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2429 = {{7'd0}, _T_14417}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14460 = _T_14458 + _GEN_2429; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_118; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2432 = {{1{spriteYPositionReg_118[9]}},spriteYPositionReg_118}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14486; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_118 = _T_14486[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14510 = {{1{inSpriteY_118[10]}},inSpriteY_118}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14528 = inSpriteX_118; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14536 = {{2'd0}, _T_14528}; // @[Mux.scala 80:57]
  wire [11:0] _T_14540 = {{1{inSpriteY_118[10]}},inSpriteY_118}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14548 = {{2'd0}, _T_14540}; // @[Mux.scala 80:57]
  wire  _T_14549 = $signed(inSpriteX_118) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14550 = $signed(inSpriteX_118) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14551 = _T_14549 & _T_14550; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14552 = $signed(_T_14510) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14553 = $signed(_T_14510) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14554 = _T_14552 & _T_14553; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14577 = _T_14548 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2438 = {{7'd0}, _T_14536}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14579 = _T_14577 + _GEN_2438; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_119; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2441 = {{1{spriteYPositionReg_119[9]}},spriteYPositionReg_119}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14605; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_119 = _T_14605[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14629 = {{1{inSpriteY_119[10]}},inSpriteY_119}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14647 = inSpriteX_119; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14655 = {{2'd0}, _T_14647}; // @[Mux.scala 80:57]
  wire [11:0] _T_14659 = {{1{inSpriteY_119[10]}},inSpriteY_119}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14667 = {{2'd0}, _T_14659}; // @[Mux.scala 80:57]
  wire  _T_14668 = $signed(inSpriteX_119) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14669 = $signed(inSpriteX_119) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14670 = _T_14668 & _T_14669; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14671 = $signed(_T_14629) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14672 = $signed(_T_14629) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14673 = _T_14671 & _T_14672; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14696 = _T_14667 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2447 = {{7'd0}, _T_14655}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14698 = _T_14696 + _GEN_2447; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_120; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2450 = {{1{spriteYPositionReg_120[9]}},spriteYPositionReg_120}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14724; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_120 = _T_14724[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14748 = {{1{inSpriteY_120[10]}},inSpriteY_120}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14766 = inSpriteX_120; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14774 = {{2'd0}, _T_14766}; // @[Mux.scala 80:57]
  wire [11:0] _T_14778 = {{1{inSpriteY_120[10]}},inSpriteY_120}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14786 = {{2'd0}, _T_14778}; // @[Mux.scala 80:57]
  wire  _T_14787 = $signed(inSpriteX_120) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14788 = $signed(inSpriteX_120) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14789 = _T_14787 & _T_14788; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14790 = $signed(_T_14748) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14791 = $signed(_T_14748) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14792 = _T_14790 & _T_14791; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14815 = _T_14786 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2456 = {{7'd0}, _T_14774}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14817 = _T_14815 + _GEN_2456; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_121; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2459 = {{1{spriteYPositionReg_121[9]}},spriteYPositionReg_121}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14843; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_121 = _T_14843[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14867 = {{1{inSpriteY_121[10]}},inSpriteY_121}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14885 = inSpriteX_121; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_14893 = {{2'd0}, _T_14885}; // @[Mux.scala 80:57]
  wire [11:0] _T_14897 = {{1{inSpriteY_121[10]}},inSpriteY_121}; // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_14905 = {{2'd0}, _T_14897}; // @[Mux.scala 80:57]
  wire  _T_14906 = $signed(inSpriteX_121) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_14907 = $signed(inSpriteX_121) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_14908 = _T_14906 & _T_14907; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_14909 = $signed(_T_14867) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_14910 = $signed(_T_14867) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_14911 = _T_14909 & _T_14910; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_14934 = _T_14905 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2465 = {{7'd0}, _T_14893}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_14936 = _T_14934 + _GEN_2465; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_122; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2468 = {{1{spriteYPositionReg_122[9]}},spriteYPositionReg_122}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_14962; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_122 = _T_14962[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_14986 = {{1{inSpriteY_122[10]}},inSpriteY_122}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_14999 = $signed(_GEN_1378) - $signed(_T_14986); // @[GraphicEngineVGA.scala 373:65]
  wire [11:0] _T_15000 = spriteFlipVerticalReg_122 ? $signed(_T_14999) : $signed(_T_14986); // @[GraphicEngineVGA.scala 373:23]
  wire [11:0] _T_15004 = inSpriteX_122; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_15012 = {{2'd0}, _T_15004}; // @[Mux.scala 80:57]
  wire [11:0] _T_15016 = spriteFlipVerticalReg_122 ? $signed(_T_14999) : $signed(_T_14986); // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_15024 = {{2'd0}, _T_15016}; // @[Mux.scala 80:57]
  wire  _T_15025 = $signed(inSpriteX_122) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_15026 = $signed(inSpriteX_122) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_15027 = _T_15025 & _T_15026; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_15028 = $signed(_T_15000) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_15029 = $signed(_T_15000) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_15030 = _T_15028 & _T_15029; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_15053 = _T_15024 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2474 = {{7'd0}, _T_15012}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_15055 = _T_15053 + _GEN_2474; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_123; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2477 = {{1{spriteYPositionReg_123[9]}},spriteYPositionReg_123}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_15081; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_123 = _T_15081[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_15105 = {{1{inSpriteY_123[10]}},inSpriteY_123}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_15118 = $signed(_GEN_1378) - $signed(_T_15105); // @[GraphicEngineVGA.scala 373:65]
  wire [11:0] _T_15119 = spriteFlipVerticalReg_123 ? $signed(_T_15118) : $signed(_T_15105); // @[GraphicEngineVGA.scala 373:23]
  wire [11:0] _T_15123 = inSpriteX_123; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_15131 = {{2'd0}, _T_15123}; // @[Mux.scala 80:57]
  wire [11:0] _T_15135 = spriteFlipVerticalReg_123 ? $signed(_T_15118) : $signed(_T_15105); // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_15143 = {{2'd0}, _T_15135}; // @[Mux.scala 80:57]
  wire  _T_15144 = $signed(inSpriteX_123) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_15145 = $signed(inSpriteX_123) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_15146 = _T_15144 & _T_15145; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_15147 = $signed(_T_15119) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_15148 = $signed(_T_15119) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_15149 = _T_15147 & _T_15148; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_15172 = _T_15143 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2483 = {{7'd0}, _T_15131}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_15174 = _T_15172 + _GEN_2483; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_124; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2486 = {{1{spriteYPositionReg_124[9]}},spriteYPositionReg_124}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_15200; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_124 = _T_15200[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_15224 = {{1{inSpriteY_124[10]}},inSpriteY_124}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_15237 = $signed(_GEN_1378) - $signed(_T_15224); // @[GraphicEngineVGA.scala 373:65]
  wire [11:0] _T_15238 = spriteFlipVerticalReg_124 ? $signed(_T_15237) : $signed(_T_15224); // @[GraphicEngineVGA.scala 373:23]
  wire [11:0] _T_15242 = inSpriteX_124; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_15250 = {{2'd0}, _T_15242}; // @[Mux.scala 80:57]
  wire [11:0] _T_15254 = spriteFlipVerticalReg_124 ? $signed(_T_15237) : $signed(_T_15224); // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_15262 = {{2'd0}, _T_15254}; // @[Mux.scala 80:57]
  wire  _T_15263 = $signed(inSpriteX_124) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_15264 = $signed(inSpriteX_124) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_15265 = _T_15263 & _T_15264; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_15266 = $signed(_T_15238) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_15267 = $signed(_T_15238) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_15268 = _T_15266 & _T_15267; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_15291 = _T_15262 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2492 = {{7'd0}, _T_15250}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_15293 = _T_15291 + _GEN_2492; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_125; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2495 = {{1{spriteYPositionReg_125[9]}},spriteYPositionReg_125}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_15319; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_125 = _T_15319[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_15343 = {{1{inSpriteY_125[10]}},inSpriteY_125}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_15356 = $signed(_GEN_1378) - $signed(_T_15343); // @[GraphicEngineVGA.scala 373:65]
  wire [11:0] _T_15357 = spriteFlipVerticalReg_125 ? $signed(_T_15356) : $signed(_T_15343); // @[GraphicEngineVGA.scala 373:23]
  wire [11:0] _T_15361 = inSpriteX_125; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_15369 = {{2'd0}, _T_15361}; // @[Mux.scala 80:57]
  wire [11:0] _T_15373 = spriteFlipVerticalReg_125 ? $signed(_T_15356) : $signed(_T_15343); // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_15381 = {{2'd0}, _T_15373}; // @[Mux.scala 80:57]
  wire  _T_15382 = $signed(inSpriteX_125) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_15383 = $signed(inSpriteX_125) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_15384 = _T_15382 & _T_15383; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_15385 = $signed(_T_15357) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_15386 = $signed(_T_15357) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_15387 = _T_15385 & _T_15386; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_15410 = _T_15381 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2501 = {{7'd0}, _T_15369}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_15412 = _T_15410 + _GEN_2501; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_126; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2504 = {{1{spriteYPositionReg_126[9]}},spriteYPositionReg_126}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_15438; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_126 = _T_15438[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_15462 = {{1{inSpriteY_126[10]}},inSpriteY_126}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_15475 = $signed(_GEN_1378) - $signed(_T_15462); // @[GraphicEngineVGA.scala 373:65]
  wire [11:0] _T_15476 = spriteFlipVerticalReg_126 ? $signed(_T_15475) : $signed(_T_15462); // @[GraphicEngineVGA.scala 373:23]
  wire [11:0] _T_15480 = inSpriteX_126; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_15488 = {{2'd0}, _T_15480}; // @[Mux.scala 80:57]
  wire [11:0] _T_15492 = spriteFlipVerticalReg_126 ? $signed(_T_15475) : $signed(_T_15462); // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_15500 = {{2'd0}, _T_15492}; // @[Mux.scala 80:57]
  wire  _T_15501 = $signed(inSpriteX_126) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_15502 = $signed(inSpriteX_126) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_15503 = _T_15501 & _T_15502; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_15504 = $signed(_T_15476) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_15505 = $signed(_T_15476) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_15506 = _T_15504 & _T_15505; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_15529 = _T_15500 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2510 = {{7'd0}, _T_15488}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_15531 = _T_15529 + _GEN_2510; // @[GraphicEngineVGA.scala 399:51]
  reg [11:0] inSpriteX_127; // @[GraphicEngineVGA.scala 355:30]
  wire [10:0] _GEN_2513 = {{1{spriteYPositionReg_127[9]}},spriteYPositionReg_127}; // @[GraphicEngineVGA.scala 356:59]
  reg [11:0] _T_15557; // @[GraphicEngineVGA.scala 356:30]
  wire [10:0] inSpriteY_127 = _T_15557[10:0]; // @[GraphicEngineVGA.scala 330:23 GraphicEngineVGA.scala 356:20]
  wire [11:0] _T_15581 = {{1{inSpriteY_127[10]}},inSpriteY_127}; // @[GraphicEngineVGA.scala 370:21]
  wire [11:0] _T_15594 = $signed(_GEN_1378) - $signed(_T_15581); // @[GraphicEngineVGA.scala 373:65]
  wire [11:0] _T_15595 = spriteFlipVerticalReg_127 ? $signed(_T_15594) : $signed(_T_15581); // @[GraphicEngineVGA.scala 373:23]
  wire [11:0] _T_15599 = inSpriteX_127; // @[GraphicEngineVGA.scala 380:24]
  wire [13:0] _T_15607 = {{2'd0}, _T_15599}; // @[Mux.scala 80:57]
  wire [11:0] _T_15611 = spriteFlipVerticalReg_127 ? $signed(_T_15594) : $signed(_T_15581); // @[GraphicEngineVGA.scala 386:24]
  wire [13:0] _T_15619 = {{2'd0}, _T_15611}; // @[Mux.scala 80:57]
  wire  _T_15620 = $signed(inSpriteX_127) >= 12'sh0; // @[GraphicEngineVGA.scala 391:31]
  wire  _T_15621 = $signed(inSpriteX_127) < 12'sh20; // @[GraphicEngineVGA.scala 391:52]
  wire  _T_15622 = _T_15620 & _T_15621; // @[GraphicEngineVGA.scala 391:39]
  wire  _T_15623 = $signed(_T_15595) >= 12'sh0; // @[GraphicEngineVGA.scala 392:31]
  wire  _T_15624 = $signed(_T_15595) < 12'sh20; // @[GraphicEngineVGA.scala 392:52]
  wire  _T_15625 = _T_15623 & _T_15624; // @[GraphicEngineVGA.scala 392:39]
  wire [20:0] _T_15648 = _T_15619 * 14'h20; // @[GraphicEngineVGA.scala 399:27]
  wire [20:0] _GEN_2519 = {{7'd0}, _T_15607}; // @[GraphicEngineVGA.scala 399:51]
  wire [20:0] _T_15650 = _T_15648 + _GEN_2519; // @[GraphicEngineVGA.scala 399:51]
  reg  _T_15660_0; // @[GameUtilities.scala 21:24]
  reg  _T_15660_1; // @[GameUtilities.scala 21:24]
  reg  _T_15660_2; // @[GameUtilities.scala 21:24]
  reg  _T_15662_0; // @[GameUtilities.scala 21:24]
  reg  _T_15662_1; // @[GameUtilities.scala 21:24]
  reg  _T_15662_2; // @[GameUtilities.scala 21:24]
  reg  _T_15664_0; // @[GameUtilities.scala 21:24]
  reg  _T_15664_1; // @[GameUtilities.scala 21:24]
  reg  _T_15664_2; // @[GameUtilities.scala 21:24]
  Memory backTileMemories_0_0 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_0_clock),
    .io_address(backTileMemories_0_0_io_address),
    .io_dataRead(backTileMemories_0_0_io_dataRead)
  );
  Memory_1 backTileMemories_0_1 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_1_clock),
    .io_address(backTileMemories_0_1_io_address),
    .io_dataRead(backTileMemories_0_1_io_dataRead)
  );
  Memory_2 backTileMemories_0_2 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_2_clock),
    .io_address(backTileMemories_0_2_io_address),
    .io_dataRead(backTileMemories_0_2_io_dataRead)
  );
  Memory_3 backTileMemories_0_3 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_3_clock),
    .io_address(backTileMemories_0_3_io_address),
    .io_dataRead(backTileMemories_0_3_io_dataRead)
  );
  Memory_4 backTileMemories_0_4 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_4_clock),
    .io_address(backTileMemories_0_4_io_address),
    .io_dataRead(backTileMemories_0_4_io_dataRead)
  );
  Memory_5 backTileMemories_0_5 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_5_clock),
    .io_address(backTileMemories_0_5_io_address),
    .io_dataRead(backTileMemories_0_5_io_dataRead)
  );
  Memory_6 backTileMemories_0_6 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_6_clock),
    .io_address(backTileMemories_0_6_io_address),
    .io_dataRead(backTileMemories_0_6_io_dataRead)
  );
  Memory_7 backTileMemories_0_7 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_7_clock),
    .io_address(backTileMemories_0_7_io_address),
    .io_dataRead(backTileMemories_0_7_io_dataRead)
  );
  Memory_8 backTileMemories_0_8 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_8_clock),
    .io_address(backTileMemories_0_8_io_address),
    .io_dataRead(backTileMemories_0_8_io_dataRead)
  );
  Memory_9 backTileMemories_0_9 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_9_clock),
    .io_address(backTileMemories_0_9_io_address),
    .io_dataRead(backTileMemories_0_9_io_dataRead)
  );
  Memory_10 backTileMemories_0_10 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_10_clock),
    .io_address(backTileMemories_0_10_io_address),
    .io_dataRead(backTileMemories_0_10_io_dataRead)
  );
  Memory_11 backTileMemories_0_11 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_11_clock),
    .io_address(backTileMemories_0_11_io_address),
    .io_dataRead(backTileMemories_0_11_io_dataRead)
  );
  Memory_12 backTileMemories_0_12 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_12_clock),
    .io_address(backTileMemories_0_12_io_address),
    .io_dataRead(backTileMemories_0_12_io_dataRead)
  );
  Memory_13 backTileMemories_0_13 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_13_clock),
    .io_address(backTileMemories_0_13_io_address),
    .io_dataRead(backTileMemories_0_13_io_dataRead)
  );
  Memory_14 backTileMemories_0_14 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_14_clock),
    .io_address(backTileMemories_0_14_io_address),
    .io_dataRead(backTileMemories_0_14_io_dataRead)
  );
  Memory_15 backTileMemories_0_15 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_15_clock),
    .io_address(backTileMemories_0_15_io_address),
    .io_dataRead(backTileMemories_0_15_io_dataRead)
  );
  Memory_16 backTileMemories_0_16 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_16_clock),
    .io_address(backTileMemories_0_16_io_address),
    .io_dataRead(backTileMemories_0_16_io_dataRead)
  );
  Memory_17 backTileMemories_0_17 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_17_clock),
    .io_address(backTileMemories_0_17_io_address),
    .io_dataRead(backTileMemories_0_17_io_dataRead)
  );
  Memory_18 backTileMemories_0_18 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_18_clock),
    .io_address(backTileMemories_0_18_io_address),
    .io_dataRead(backTileMemories_0_18_io_dataRead)
  );
  Memory_19 backTileMemories_0_19 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_19_clock),
    .io_address(backTileMemories_0_19_io_address),
    .io_dataRead(backTileMemories_0_19_io_dataRead)
  );
  Memory_20 backTileMemories_0_20 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_20_clock),
    .io_address(backTileMemories_0_20_io_address),
    .io_dataRead(backTileMemories_0_20_io_dataRead)
  );
  Memory_21 backTileMemories_0_21 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_21_clock),
    .io_address(backTileMemories_0_21_io_address),
    .io_dataRead(backTileMemories_0_21_io_dataRead)
  );
  Memory_22 backTileMemories_0_22 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_22_clock),
    .io_address(backTileMemories_0_22_io_address),
    .io_dataRead(backTileMemories_0_22_io_dataRead)
  );
  Memory_23 backTileMemories_0_23 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_23_clock),
    .io_address(backTileMemories_0_23_io_address),
    .io_dataRead(backTileMemories_0_23_io_dataRead)
  );
  Memory_24 backTileMemories_0_24 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_24_clock),
    .io_address(backTileMemories_0_24_io_address),
    .io_dataRead(backTileMemories_0_24_io_dataRead)
  );
  Memory_25 backTileMemories_0_25 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_25_clock),
    .io_address(backTileMemories_0_25_io_address),
    .io_dataRead(backTileMemories_0_25_io_dataRead)
  );
  Memory_26 backTileMemories_0_26 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_26_clock),
    .io_address(backTileMemories_0_26_io_address),
    .io_dataRead(backTileMemories_0_26_io_dataRead)
  );
  Memory_27 backTileMemories_0_27 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_27_clock),
    .io_address(backTileMemories_0_27_io_address),
    .io_dataRead(backTileMemories_0_27_io_dataRead)
  );
  Memory_28 backTileMemories_0_28 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_28_clock),
    .io_address(backTileMemories_0_28_io_address),
    .io_dataRead(backTileMemories_0_28_io_dataRead)
  );
  Memory_29 backTileMemories_0_29 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_29_clock),
    .io_address(backTileMemories_0_29_io_address),
    .io_dataRead(backTileMemories_0_29_io_dataRead)
  );
  Memory_30 backTileMemories_0_30 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_30_clock),
    .io_address(backTileMemories_0_30_io_address),
    .io_dataRead(backTileMemories_0_30_io_dataRead)
  );
  Memory_31 backTileMemories_0_31 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_0_31_clock),
    .io_address(backTileMemories_0_31_io_address),
    .io_dataRead(backTileMemories_0_31_io_dataRead)
  );
  Memory backTileMemories_1_0 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_0_clock),
    .io_address(backTileMemories_1_0_io_address),
    .io_dataRead(backTileMemories_1_0_io_dataRead)
  );
  Memory_1 backTileMemories_1_1 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_1_clock),
    .io_address(backTileMemories_1_1_io_address),
    .io_dataRead(backTileMemories_1_1_io_dataRead)
  );
  Memory_2 backTileMemories_1_2 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_2_clock),
    .io_address(backTileMemories_1_2_io_address),
    .io_dataRead(backTileMemories_1_2_io_dataRead)
  );
  Memory_3 backTileMemories_1_3 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_3_clock),
    .io_address(backTileMemories_1_3_io_address),
    .io_dataRead(backTileMemories_1_3_io_dataRead)
  );
  Memory_4 backTileMemories_1_4 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_4_clock),
    .io_address(backTileMemories_1_4_io_address),
    .io_dataRead(backTileMemories_1_4_io_dataRead)
  );
  Memory_5 backTileMemories_1_5 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_5_clock),
    .io_address(backTileMemories_1_5_io_address),
    .io_dataRead(backTileMemories_1_5_io_dataRead)
  );
  Memory_6 backTileMemories_1_6 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_6_clock),
    .io_address(backTileMemories_1_6_io_address),
    .io_dataRead(backTileMemories_1_6_io_dataRead)
  );
  Memory_7 backTileMemories_1_7 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_7_clock),
    .io_address(backTileMemories_1_7_io_address),
    .io_dataRead(backTileMemories_1_7_io_dataRead)
  );
  Memory_8 backTileMemories_1_8 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_8_clock),
    .io_address(backTileMemories_1_8_io_address),
    .io_dataRead(backTileMemories_1_8_io_dataRead)
  );
  Memory_9 backTileMemories_1_9 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_9_clock),
    .io_address(backTileMemories_1_9_io_address),
    .io_dataRead(backTileMemories_1_9_io_dataRead)
  );
  Memory_10 backTileMemories_1_10 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_10_clock),
    .io_address(backTileMemories_1_10_io_address),
    .io_dataRead(backTileMemories_1_10_io_dataRead)
  );
  Memory_11 backTileMemories_1_11 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_11_clock),
    .io_address(backTileMemories_1_11_io_address),
    .io_dataRead(backTileMemories_1_11_io_dataRead)
  );
  Memory_12 backTileMemories_1_12 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_12_clock),
    .io_address(backTileMemories_1_12_io_address),
    .io_dataRead(backTileMemories_1_12_io_dataRead)
  );
  Memory_13 backTileMemories_1_13 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_13_clock),
    .io_address(backTileMemories_1_13_io_address),
    .io_dataRead(backTileMemories_1_13_io_dataRead)
  );
  Memory_14 backTileMemories_1_14 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_14_clock),
    .io_address(backTileMemories_1_14_io_address),
    .io_dataRead(backTileMemories_1_14_io_dataRead)
  );
  Memory_15 backTileMemories_1_15 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_15_clock),
    .io_address(backTileMemories_1_15_io_address),
    .io_dataRead(backTileMemories_1_15_io_dataRead)
  );
  Memory_16 backTileMemories_1_16 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_16_clock),
    .io_address(backTileMemories_1_16_io_address),
    .io_dataRead(backTileMemories_1_16_io_dataRead)
  );
  Memory_17 backTileMemories_1_17 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_17_clock),
    .io_address(backTileMemories_1_17_io_address),
    .io_dataRead(backTileMemories_1_17_io_dataRead)
  );
  Memory_18 backTileMemories_1_18 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_18_clock),
    .io_address(backTileMemories_1_18_io_address),
    .io_dataRead(backTileMemories_1_18_io_dataRead)
  );
  Memory_19 backTileMemories_1_19 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_19_clock),
    .io_address(backTileMemories_1_19_io_address),
    .io_dataRead(backTileMemories_1_19_io_dataRead)
  );
  Memory_20 backTileMemories_1_20 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_20_clock),
    .io_address(backTileMemories_1_20_io_address),
    .io_dataRead(backTileMemories_1_20_io_dataRead)
  );
  Memory_21 backTileMemories_1_21 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_21_clock),
    .io_address(backTileMemories_1_21_io_address),
    .io_dataRead(backTileMemories_1_21_io_dataRead)
  );
  Memory_22 backTileMemories_1_22 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_22_clock),
    .io_address(backTileMemories_1_22_io_address),
    .io_dataRead(backTileMemories_1_22_io_dataRead)
  );
  Memory_23 backTileMemories_1_23 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_23_clock),
    .io_address(backTileMemories_1_23_io_address),
    .io_dataRead(backTileMemories_1_23_io_dataRead)
  );
  Memory_24 backTileMemories_1_24 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_24_clock),
    .io_address(backTileMemories_1_24_io_address),
    .io_dataRead(backTileMemories_1_24_io_dataRead)
  );
  Memory_25 backTileMemories_1_25 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_25_clock),
    .io_address(backTileMemories_1_25_io_address),
    .io_dataRead(backTileMemories_1_25_io_dataRead)
  );
  Memory_26 backTileMemories_1_26 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_26_clock),
    .io_address(backTileMemories_1_26_io_address),
    .io_dataRead(backTileMemories_1_26_io_dataRead)
  );
  Memory_27 backTileMemories_1_27 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_27_clock),
    .io_address(backTileMemories_1_27_io_address),
    .io_dataRead(backTileMemories_1_27_io_dataRead)
  );
  Memory_28 backTileMemories_1_28 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_28_clock),
    .io_address(backTileMemories_1_28_io_address),
    .io_dataRead(backTileMemories_1_28_io_dataRead)
  );
  Memory_29 backTileMemories_1_29 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_29_clock),
    .io_address(backTileMemories_1_29_io_address),
    .io_dataRead(backTileMemories_1_29_io_dataRead)
  );
  Memory_30 backTileMemories_1_30 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_30_clock),
    .io_address(backTileMemories_1_30_io_address),
    .io_dataRead(backTileMemories_1_30_io_dataRead)
  );
  Memory_31 backTileMemories_1_31 ( // @[GraphicEngineVGA.scala 205:34]
    .clock(backTileMemories_1_31_clock),
    .io_address(backTileMemories_1_31_io_address),
    .io_dataRead(backTileMemories_1_31_io_dataRead)
  );
  Memory_64 backBufferMemories_0 ( // @[GraphicEngineVGA.scala 230:34]
    .clock(backBufferMemories_0_clock),
    .io_address(backBufferMemories_0_io_address),
    .io_dataRead(backBufferMemories_0_io_dataRead),
    .io_writeEnable(backBufferMemories_0_io_writeEnable),
    .io_dataWrite(backBufferMemories_0_io_dataWrite)
  );
  Memory_64 backBufferMemories_1 ( // @[GraphicEngineVGA.scala 230:34]
    .clock(backBufferMemories_1_clock),
    .io_address(backBufferMemories_1_io_address),
    .io_dataRead(backBufferMemories_1_io_dataRead),
    .io_writeEnable(backBufferMemories_1_io_writeEnable),
    .io_dataWrite(backBufferMemories_1_io_dataWrite)
  );
  Memory_64 backBufferShadowMemories_0 ( // @[GraphicEngineVGA.scala 235:40]
    .clock(backBufferShadowMemories_0_clock),
    .io_address(backBufferShadowMemories_0_io_address),
    .io_dataRead(backBufferShadowMemories_0_io_dataRead),
    .io_writeEnable(backBufferShadowMemories_0_io_writeEnable),
    .io_dataWrite(backBufferShadowMemories_0_io_dataWrite)
  );
  Memory_64 backBufferShadowMemories_1 ( // @[GraphicEngineVGA.scala 235:40]
    .clock(backBufferShadowMemories_1_clock),
    .io_address(backBufferShadowMemories_1_io_address),
    .io_dataRead(backBufferShadowMemories_1_io_dataRead),
    .io_writeEnable(backBufferShadowMemories_1_io_writeEnable),
    .io_dataWrite(backBufferShadowMemories_1_io_dataWrite)
  );
  Memory_68 backBufferRestoreMemories_0 ( // @[GraphicEngineVGA.scala 241:41]
    .clock(backBufferRestoreMemories_0_clock),
    .io_address(backBufferRestoreMemories_0_io_address),
    .io_dataRead(backBufferRestoreMemories_0_io_dataRead)
  );
  Memory_69 backBufferRestoreMemories_1 ( // @[GraphicEngineVGA.scala 241:41]
    .clock(backBufferRestoreMemories_1_clock),
    .io_address(backBufferRestoreMemories_1_io_address),
    .io_dataRead(backBufferRestoreMemories_1_io_dataRead)
  );
  Memory_70 spriteMemories_0 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_0_clock),
    .io_address(spriteMemories_0_io_address),
    .io_dataRead(spriteMemories_0_io_dataRead)
  );
  Memory_71 spriteMemories_1 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_1_clock),
    .io_address(spriteMemories_1_io_address),
    .io_dataRead(spriteMemories_1_io_dataRead)
  );
  Memory_72 spriteMemories_2 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_2_clock),
    .io_address(spriteMemories_2_io_address),
    .io_dataRead(spriteMemories_2_io_dataRead)
  );
  Memory_73 spriteMemories_3 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_3_clock),
    .io_address(spriteMemories_3_io_address),
    .io_dataRead(spriteMemories_3_io_dataRead)
  );
  Memory_74 spriteMemories_4 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_4_clock),
    .io_address(spriteMemories_4_io_address),
    .io_dataRead(spriteMemories_4_io_dataRead)
  );
  Memory_75 spriteMemories_5 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_5_clock),
    .io_address(spriteMemories_5_io_address),
    .io_dataRead(spriteMemories_5_io_dataRead)
  );
  Memory_76 spriteMemories_6 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_6_clock),
    .io_address(spriteMemories_6_io_address),
    .io_dataRead(spriteMemories_6_io_dataRead)
  );
  Memory_77 spriteMemories_7 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_7_clock),
    .io_address(spriteMemories_7_io_address),
    .io_dataRead(spriteMemories_7_io_dataRead)
  );
  Memory_78 spriteMemories_8 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_8_clock),
    .io_address(spriteMemories_8_io_address),
    .io_dataRead(spriteMemories_8_io_dataRead)
  );
  Memory_79 spriteMemories_9 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_9_clock),
    .io_address(spriteMemories_9_io_address),
    .io_dataRead(spriteMemories_9_io_dataRead)
  );
  Memory_80 spriteMemories_10 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_10_clock),
    .io_address(spriteMemories_10_io_address),
    .io_dataRead(spriteMemories_10_io_dataRead)
  );
  Memory_81 spriteMemories_11 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_11_clock),
    .io_address(spriteMemories_11_io_address),
    .io_dataRead(spriteMemories_11_io_dataRead)
  );
  Memory_82 spriteMemories_12 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_12_clock),
    .io_address(spriteMemories_12_io_address),
    .io_dataRead(spriteMemories_12_io_dataRead)
  );
  Memory_83 spriteMemories_13 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_13_clock),
    .io_address(spriteMemories_13_io_address),
    .io_dataRead(spriteMemories_13_io_dataRead)
  );
  Memory_84 spriteMemories_14 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_14_clock),
    .io_address(spriteMemories_14_io_address),
    .io_dataRead(spriteMemories_14_io_dataRead)
  );
  Memory_85 spriteMemories_15 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_15_clock),
    .io_address(spriteMemories_15_io_address),
    .io_dataRead(spriteMemories_15_io_dataRead)
  );
  Memory_86 spriteMemories_16 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_16_clock),
    .io_address(spriteMemories_16_io_address),
    .io_dataRead(spriteMemories_16_io_dataRead)
  );
  Memory_87 spriteMemories_17 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_17_clock),
    .io_address(spriteMemories_17_io_address),
    .io_dataRead(spriteMemories_17_io_dataRead)
  );
  Memory_88 spriteMemories_18 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_18_clock),
    .io_address(spriteMemories_18_io_address),
    .io_dataRead(spriteMemories_18_io_dataRead)
  );
  Memory_89 spriteMemories_19 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_19_clock),
    .io_address(spriteMemories_19_io_address),
    .io_dataRead(spriteMemories_19_io_dataRead)
  );
  Memory_90 spriteMemories_20 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_20_clock),
    .io_address(spriteMemories_20_io_address),
    .io_dataRead(spriteMemories_20_io_dataRead)
  );
  Memory_91 spriteMemories_21 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_21_clock),
    .io_address(spriteMemories_21_io_address),
    .io_dataRead(spriteMemories_21_io_dataRead)
  );
  Memory_92 spriteMemories_22 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_22_clock),
    .io_address(spriteMemories_22_io_address),
    .io_dataRead(spriteMemories_22_io_dataRead)
  );
  Memory_93 spriteMemories_23 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_23_clock),
    .io_address(spriteMemories_23_io_address),
    .io_dataRead(spriteMemories_23_io_dataRead)
  );
  Memory_94 spriteMemories_24 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_24_clock),
    .io_address(spriteMemories_24_io_address),
    .io_dataRead(spriteMemories_24_io_dataRead)
  );
  Memory_95 spriteMemories_25 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_25_clock),
    .io_address(spriteMemories_25_io_address),
    .io_dataRead(spriteMemories_25_io_dataRead)
  );
  Memory_96 spriteMemories_26 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_26_clock),
    .io_address(spriteMemories_26_io_address),
    .io_dataRead(spriteMemories_26_io_dataRead)
  );
  Memory_97 spriteMemories_27 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_27_clock),
    .io_address(spriteMemories_27_io_address),
    .io_dataRead(spriteMemories_27_io_dataRead)
  );
  Memory_98 spriteMemories_28 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_28_clock),
    .io_address(spriteMemories_28_io_address),
    .io_dataRead(spriteMemories_28_io_dataRead)
  );
  Memory_99 spriteMemories_29 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_29_clock),
    .io_address(spriteMemories_29_io_address),
    .io_dataRead(spriteMemories_29_io_dataRead)
  );
  Memory_100 spriteMemories_30 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_30_clock),
    .io_address(spriteMemories_30_io_address),
    .io_dataRead(spriteMemories_30_io_dataRead)
  );
  Memory_101 spriteMemories_31 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_31_clock),
    .io_address(spriteMemories_31_io_address),
    .io_dataRead(spriteMemories_31_io_dataRead)
  );
  Memory_102 spriteMemories_32 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_32_clock),
    .io_address(spriteMemories_32_io_address),
    .io_dataRead(spriteMemories_32_io_dataRead)
  );
  Memory_103 spriteMemories_33 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_33_clock),
    .io_address(spriteMemories_33_io_address),
    .io_dataRead(spriteMemories_33_io_dataRead)
  );
  Memory_104 spriteMemories_34 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_34_clock),
    .io_address(spriteMemories_34_io_address),
    .io_dataRead(spriteMemories_34_io_dataRead)
  );
  Memory_105 spriteMemories_35 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_35_clock),
    .io_address(spriteMemories_35_io_address),
    .io_dataRead(spriteMemories_35_io_dataRead)
  );
  Memory_106 spriteMemories_36 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_36_clock),
    .io_address(spriteMemories_36_io_address),
    .io_dataRead(spriteMemories_36_io_dataRead)
  );
  Memory_107 spriteMemories_37 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_37_clock),
    .io_address(spriteMemories_37_io_address),
    .io_dataRead(spriteMemories_37_io_dataRead)
  );
  Memory_108 spriteMemories_38 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_38_clock),
    .io_address(spriteMemories_38_io_address),
    .io_dataRead(spriteMemories_38_io_dataRead)
  );
  Memory_109 spriteMemories_39 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_39_clock),
    .io_address(spriteMemories_39_io_address),
    .io_dataRead(spriteMemories_39_io_dataRead)
  );
  Memory_110 spriteMemories_40 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_40_clock),
    .io_address(spriteMemories_40_io_address),
    .io_dataRead(spriteMemories_40_io_dataRead)
  );
  Memory_111 spriteMemories_41 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_41_clock),
    .io_address(spriteMemories_41_io_address),
    .io_dataRead(spriteMemories_41_io_dataRead)
  );
  Memory_112 spriteMemories_42 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_42_clock),
    .io_address(spriteMemories_42_io_address),
    .io_dataRead(spriteMemories_42_io_dataRead)
  );
  Memory_113 spriteMemories_43 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_43_clock),
    .io_address(spriteMemories_43_io_address),
    .io_dataRead(spriteMemories_43_io_dataRead)
  );
  Memory_114 spriteMemories_44 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_44_clock),
    .io_address(spriteMemories_44_io_address),
    .io_dataRead(spriteMemories_44_io_dataRead)
  );
  Memory_115 spriteMemories_45 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_45_clock),
    .io_address(spriteMemories_45_io_address),
    .io_dataRead(spriteMemories_45_io_dataRead)
  );
  Memory_116 spriteMemories_46 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_46_clock),
    .io_address(spriteMemories_46_io_address),
    .io_dataRead(spriteMemories_46_io_dataRead)
  );
  Memory_117 spriteMemories_47 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_47_clock),
    .io_address(spriteMemories_47_io_address),
    .io_dataRead(spriteMemories_47_io_dataRead)
  );
  Memory_118 spriteMemories_48 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_48_clock),
    .io_address(spriteMemories_48_io_address),
    .io_dataRead(spriteMemories_48_io_dataRead)
  );
  Memory_119 spriteMemories_49 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_49_clock),
    .io_address(spriteMemories_49_io_address),
    .io_dataRead(spriteMemories_49_io_dataRead)
  );
  Memory_120 spriteMemories_50 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_50_clock),
    .io_address(spriteMemories_50_io_address),
    .io_dataRead(spriteMemories_50_io_dataRead)
  );
  Memory_121 spriteMemories_51 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_51_clock),
    .io_address(spriteMemories_51_io_address),
    .io_dataRead(spriteMemories_51_io_dataRead)
  );
  Memory_122 spriteMemories_52 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_52_clock),
    .io_address(spriteMemories_52_io_address),
    .io_dataRead(spriteMemories_52_io_dataRead)
  );
  Memory_123 spriteMemories_53 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_53_clock),
    .io_address(spriteMemories_53_io_address),
    .io_dataRead(spriteMemories_53_io_dataRead)
  );
  Memory_124 spriteMemories_54 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_54_clock),
    .io_address(spriteMemories_54_io_address),
    .io_dataRead(spriteMemories_54_io_dataRead)
  );
  Memory_125 spriteMemories_55 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_55_clock),
    .io_address(spriteMemories_55_io_address),
    .io_dataRead(spriteMemories_55_io_dataRead)
  );
  Memory_126 spriteMemories_56 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_56_clock),
    .io_address(spriteMemories_56_io_address),
    .io_dataRead(spriteMemories_56_io_dataRead)
  );
  Memory_127 spriteMemories_57 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_57_clock),
    .io_address(spriteMemories_57_io_address),
    .io_dataRead(spriteMemories_57_io_dataRead)
  );
  Memory_128 spriteMemories_58 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_58_clock),
    .io_address(spriteMemories_58_io_address),
    .io_dataRead(spriteMemories_58_io_dataRead)
  );
  Memory_129 spriteMemories_59 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_59_clock),
    .io_address(spriteMemories_59_io_address),
    .io_dataRead(spriteMemories_59_io_dataRead)
  );
  Memory_130 spriteMemories_60 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_60_clock),
    .io_address(spriteMemories_60_io_address),
    .io_dataRead(spriteMemories_60_io_dataRead)
  );
  Memory_131 spriteMemories_61 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_61_clock),
    .io_address(spriteMemories_61_io_address),
    .io_dataRead(spriteMemories_61_io_dataRead)
  );
  Memory_132 spriteMemories_62 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_62_clock),
    .io_address(spriteMemories_62_io_address),
    .io_dataRead(spriteMemories_62_io_dataRead)
  );
  Memory_133 spriteMemories_63 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_63_clock),
    .io_address(spriteMemories_63_io_address),
    .io_dataRead(spriteMemories_63_io_dataRead)
  );
  Memory_134 spriteMemories_64 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_64_clock),
    .io_address(spriteMemories_64_io_address),
    .io_dataRead(spriteMemories_64_io_dataRead)
  );
  Memory_135 spriteMemories_65 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_65_clock),
    .io_address(spriteMemories_65_io_address),
    .io_dataRead(spriteMemories_65_io_dataRead)
  );
  Memory_136 spriteMemories_66 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_66_clock),
    .io_address(spriteMemories_66_io_address),
    .io_dataRead(spriteMemories_66_io_dataRead)
  );
  Memory_137 spriteMemories_67 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_67_clock),
    .io_address(spriteMemories_67_io_address),
    .io_dataRead(spriteMemories_67_io_dataRead)
  );
  Memory_138 spriteMemories_68 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_68_clock),
    .io_address(spriteMemories_68_io_address),
    .io_dataRead(spriteMemories_68_io_dataRead)
  );
  Memory_139 spriteMemories_69 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_69_clock),
    .io_address(spriteMemories_69_io_address),
    .io_dataRead(spriteMemories_69_io_dataRead)
  );
  Memory_140 spriteMemories_70 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_70_clock),
    .io_address(spriteMemories_70_io_address),
    .io_dataRead(spriteMemories_70_io_dataRead)
  );
  Memory_141 spriteMemories_71 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_71_clock),
    .io_address(spriteMemories_71_io_address),
    .io_dataRead(spriteMemories_71_io_dataRead)
  );
  Memory_142 spriteMemories_72 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_72_clock),
    .io_address(spriteMemories_72_io_address),
    .io_dataRead(spriteMemories_72_io_dataRead)
  );
  Memory_143 spriteMemories_73 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_73_clock),
    .io_address(spriteMemories_73_io_address),
    .io_dataRead(spriteMemories_73_io_dataRead)
  );
  Memory_144 spriteMemories_74 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_74_clock),
    .io_address(spriteMemories_74_io_address),
    .io_dataRead(spriteMemories_74_io_dataRead)
  );
  Memory_145 spriteMemories_75 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_75_clock),
    .io_address(spriteMemories_75_io_address),
    .io_dataRead(spriteMemories_75_io_dataRead)
  );
  Memory_146 spriteMemories_76 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_76_clock),
    .io_address(spriteMemories_76_io_address),
    .io_dataRead(spriteMemories_76_io_dataRead)
  );
  Memory_147 spriteMemories_77 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_77_clock),
    .io_address(spriteMemories_77_io_address),
    .io_dataRead(spriteMemories_77_io_dataRead)
  );
  Memory_148 spriteMemories_78 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_78_clock),
    .io_address(spriteMemories_78_io_address),
    .io_dataRead(spriteMemories_78_io_dataRead)
  );
  Memory_149 spriteMemories_79 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_79_clock),
    .io_address(spriteMemories_79_io_address),
    .io_dataRead(spriteMemories_79_io_dataRead)
  );
  Memory_150 spriteMemories_80 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_80_clock),
    .io_address(spriteMemories_80_io_address),
    .io_dataRead(spriteMemories_80_io_dataRead)
  );
  Memory_151 spriteMemories_81 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_81_clock),
    .io_address(spriteMemories_81_io_address),
    .io_dataRead(spriteMemories_81_io_dataRead)
  );
  Memory_152 spriteMemories_82 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_82_clock),
    .io_address(spriteMemories_82_io_address),
    .io_dataRead(spriteMemories_82_io_dataRead)
  );
  Memory_153 spriteMemories_83 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_83_clock),
    .io_address(spriteMemories_83_io_address),
    .io_dataRead(spriteMemories_83_io_dataRead)
  );
  Memory_154 spriteMemories_84 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_84_clock),
    .io_address(spriteMemories_84_io_address),
    .io_dataRead(spriteMemories_84_io_dataRead)
  );
  Memory_155 spriteMemories_85 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_85_clock),
    .io_address(spriteMemories_85_io_address),
    .io_dataRead(spriteMemories_85_io_dataRead)
  );
  Memory_156 spriteMemories_86 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_86_clock),
    .io_address(spriteMemories_86_io_address),
    .io_dataRead(spriteMemories_86_io_dataRead)
  );
  Memory_157 spriteMemories_87 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_87_clock),
    .io_address(spriteMemories_87_io_address),
    .io_dataRead(spriteMemories_87_io_dataRead)
  );
  Memory_158 spriteMemories_88 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_88_clock),
    .io_address(spriteMemories_88_io_address),
    .io_dataRead(spriteMemories_88_io_dataRead)
  );
  Memory_159 spriteMemories_89 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_89_clock),
    .io_address(spriteMemories_89_io_address),
    .io_dataRead(spriteMemories_89_io_dataRead)
  );
  Memory_160 spriteMemories_90 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_90_clock),
    .io_address(spriteMemories_90_io_address),
    .io_dataRead(spriteMemories_90_io_dataRead)
  );
  Memory_161 spriteMemories_91 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_91_clock),
    .io_address(spriteMemories_91_io_address),
    .io_dataRead(spriteMemories_91_io_dataRead)
  );
  Memory_162 spriteMemories_92 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_92_clock),
    .io_address(spriteMemories_92_io_address),
    .io_dataRead(spriteMemories_92_io_dataRead)
  );
  Memory_163 spriteMemories_93 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_93_clock),
    .io_address(spriteMemories_93_io_address),
    .io_dataRead(spriteMemories_93_io_dataRead)
  );
  Memory_164 spriteMemories_94 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_94_clock),
    .io_address(spriteMemories_94_io_address),
    .io_dataRead(spriteMemories_94_io_dataRead)
  );
  Memory_165 spriteMemories_95 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_95_clock),
    .io_address(spriteMemories_95_io_address),
    .io_dataRead(spriteMemories_95_io_dataRead)
  );
  Memory_166 spriteMemories_96 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_96_clock),
    .io_address(spriteMemories_96_io_address),
    .io_dataRead(spriteMemories_96_io_dataRead)
  );
  Memory_167 spriteMemories_97 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_97_clock),
    .io_address(spriteMemories_97_io_address),
    .io_dataRead(spriteMemories_97_io_dataRead)
  );
  Memory_168 spriteMemories_98 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_98_clock),
    .io_address(spriteMemories_98_io_address),
    .io_dataRead(spriteMemories_98_io_dataRead)
  );
  Memory_169 spriteMemories_99 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_99_clock),
    .io_address(spriteMemories_99_io_address),
    .io_dataRead(spriteMemories_99_io_dataRead)
  );
  Memory_170 spriteMemories_100 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_100_clock),
    .io_address(spriteMemories_100_io_address),
    .io_dataRead(spriteMemories_100_io_dataRead)
  );
  Memory_171 spriteMemories_101 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_101_clock),
    .io_address(spriteMemories_101_io_address),
    .io_dataRead(spriteMemories_101_io_dataRead)
  );
  Memory_172 spriteMemories_102 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_102_clock),
    .io_address(spriteMemories_102_io_address),
    .io_dataRead(spriteMemories_102_io_dataRead)
  );
  Memory_173 spriteMemories_103 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_103_clock),
    .io_address(spriteMemories_103_io_address),
    .io_dataRead(spriteMemories_103_io_dataRead)
  );
  Memory_174 spriteMemories_104 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_104_clock),
    .io_address(spriteMemories_104_io_address),
    .io_dataRead(spriteMemories_104_io_dataRead)
  );
  Memory_175 spriteMemories_105 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_105_clock),
    .io_address(spriteMemories_105_io_address),
    .io_dataRead(spriteMemories_105_io_dataRead)
  );
  Memory_176 spriteMemories_106 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_106_clock),
    .io_address(spriteMemories_106_io_address),
    .io_dataRead(spriteMemories_106_io_dataRead)
  );
  Memory_177 spriteMemories_107 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_107_clock),
    .io_address(spriteMemories_107_io_address),
    .io_dataRead(spriteMemories_107_io_dataRead)
  );
  Memory_178 spriteMemories_108 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_108_clock),
    .io_address(spriteMemories_108_io_address),
    .io_dataRead(spriteMemories_108_io_dataRead)
  );
  Memory_179 spriteMemories_109 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_109_clock),
    .io_address(spriteMemories_109_io_address),
    .io_dataRead(spriteMemories_109_io_dataRead)
  );
  Memory_180 spriteMemories_110 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_110_clock),
    .io_address(spriteMemories_110_io_address),
    .io_dataRead(spriteMemories_110_io_dataRead)
  );
  Memory_181 spriteMemories_111 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_111_clock),
    .io_address(spriteMemories_111_io_address),
    .io_dataRead(spriteMemories_111_io_dataRead)
  );
  Memory_182 spriteMemories_112 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_112_clock),
    .io_address(spriteMemories_112_io_address),
    .io_dataRead(spriteMemories_112_io_dataRead)
  );
  Memory_183 spriteMemories_113 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_113_clock),
    .io_address(spriteMemories_113_io_address),
    .io_dataRead(spriteMemories_113_io_dataRead)
  );
  Memory_184 spriteMemories_114 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_114_clock),
    .io_address(spriteMemories_114_io_address),
    .io_dataRead(spriteMemories_114_io_dataRead)
  );
  Memory_185 spriteMemories_115 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_115_clock),
    .io_address(spriteMemories_115_io_address),
    .io_dataRead(spriteMemories_115_io_dataRead)
  );
  Memory_186 spriteMemories_116 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_116_clock),
    .io_address(spriteMemories_116_io_address),
    .io_dataRead(spriteMemories_116_io_dataRead)
  );
  Memory_187 spriteMemories_117 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_117_clock),
    .io_address(spriteMemories_117_io_address),
    .io_dataRead(spriteMemories_117_io_dataRead)
  );
  Memory_188 spriteMemories_118 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_118_clock),
    .io_address(spriteMemories_118_io_address),
    .io_dataRead(spriteMemories_118_io_dataRead)
  );
  Memory_189 spriteMemories_119 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_119_clock),
    .io_address(spriteMemories_119_io_address),
    .io_dataRead(spriteMemories_119_io_dataRead)
  );
  Memory_190 spriteMemories_120 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_120_clock),
    .io_address(spriteMemories_120_io_address),
    .io_dataRead(spriteMemories_120_io_dataRead)
  );
  Memory_191 spriteMemories_121 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_121_clock),
    .io_address(spriteMemories_121_io_address),
    .io_dataRead(spriteMemories_121_io_dataRead)
  );
  Memory_192 spriteMemories_122 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_122_clock),
    .io_address(spriteMemories_122_io_address),
    .io_dataRead(spriteMemories_122_io_dataRead)
  );
  Memory_193 spriteMemories_123 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_123_clock),
    .io_address(spriteMemories_123_io_address),
    .io_dataRead(spriteMemories_123_io_dataRead)
  );
  Memory_194 spriteMemories_124 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_124_clock),
    .io_address(spriteMemories_124_io_address),
    .io_dataRead(spriteMemories_124_io_dataRead)
  );
  Memory_195 spriteMemories_125 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_125_clock),
    .io_address(spriteMemories_125_io_address),
    .io_dataRead(spriteMemories_125_io_dataRead)
  );
  Memory_196 spriteMemories_126 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_126_clock),
    .io_address(spriteMemories_126_io_address),
    .io_dataRead(spriteMemories_126_io_dataRead)
  );
  Memory_197 spriteMemories_127 ( // @[GraphicEngineVGA.scala 320:30]
    .clock(spriteMemories_127_clock),
    .io_address(spriteMemories_127_io_address),
    .io_dataRead(spriteMemories_127_io_dataRead)
  );
  Memory_198 rotation45deg_0 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_0_clock),
    .io_address(rotation45deg_0_io_address)
  );
  Memory_198 rotation45deg_1 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_1_clock),
    .io_address(rotation45deg_1_io_address)
  );
  Memory_198 rotation45deg_2 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_2_clock),
    .io_address(rotation45deg_2_io_address)
  );
  Memory_198 rotation45deg_3 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_3_clock),
    .io_address(rotation45deg_3_io_address)
  );
  Memory_198 rotation45deg_4 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_4_clock),
    .io_address(rotation45deg_4_io_address)
  );
  Memory_198 rotation45deg_5 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_5_clock),
    .io_address(rotation45deg_5_io_address)
  );
  Memory_198 rotation45deg_6 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_6_clock),
    .io_address(rotation45deg_6_io_address)
  );
  Memory_198 rotation45deg_7 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_7_clock),
    .io_address(rotation45deg_7_io_address)
  );
  Memory_198 rotation45deg_8 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_8_clock),
    .io_address(rotation45deg_8_io_address)
  );
  Memory_198 rotation45deg_9 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_9_clock),
    .io_address(rotation45deg_9_io_address)
  );
  Memory_198 rotation45deg_10 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_10_clock),
    .io_address(rotation45deg_10_io_address)
  );
  Memory_198 rotation45deg_11 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_11_clock),
    .io_address(rotation45deg_11_io_address)
  );
  Memory_198 rotation45deg_12 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_12_clock),
    .io_address(rotation45deg_12_io_address)
  );
  Memory_198 rotation45deg_13 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_13_clock),
    .io_address(rotation45deg_13_io_address)
  );
  Memory_198 rotation45deg_14 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_14_clock),
    .io_address(rotation45deg_14_io_address)
  );
  Memory_198 rotation45deg_15 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_15_clock),
    .io_address(rotation45deg_15_io_address)
  );
  Memory_198 rotation45deg_16 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_16_clock),
    .io_address(rotation45deg_16_io_address)
  );
  Memory_198 rotation45deg_17 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_17_clock),
    .io_address(rotation45deg_17_io_address)
  );
  Memory_198 rotation45deg_18 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_18_clock),
    .io_address(rotation45deg_18_io_address)
  );
  Memory_198 rotation45deg_19 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_19_clock),
    .io_address(rotation45deg_19_io_address)
  );
  Memory_198 rotation45deg_20 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_20_clock),
    .io_address(rotation45deg_20_io_address)
  );
  Memory_198 rotation45deg_21 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_21_clock),
    .io_address(rotation45deg_21_io_address)
  );
  Memory_198 rotation45deg_22 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_22_clock),
    .io_address(rotation45deg_22_io_address)
  );
  Memory_198 rotation45deg_23 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_23_clock),
    .io_address(rotation45deg_23_io_address)
  );
  Memory_198 rotation45deg_24 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_24_clock),
    .io_address(rotation45deg_24_io_address)
  );
  Memory_198 rotation45deg_25 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_25_clock),
    .io_address(rotation45deg_25_io_address)
  );
  Memory_198 rotation45deg_26 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_26_clock),
    .io_address(rotation45deg_26_io_address)
  );
  Memory_198 rotation45deg_27 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_27_clock),
    .io_address(rotation45deg_27_io_address)
  );
  Memory_198 rotation45deg_28 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_28_clock),
    .io_address(rotation45deg_28_io_address)
  );
  Memory_198 rotation45deg_29 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_29_clock),
    .io_address(rotation45deg_29_io_address)
  );
  Memory_198 rotation45deg_30 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_30_clock),
    .io_address(rotation45deg_30_io_address)
  );
  Memory_198 rotation45deg_31 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_31_clock),
    .io_address(rotation45deg_31_io_address)
  );
  Memory_198 rotation45deg_32 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_32_clock),
    .io_address(rotation45deg_32_io_address)
  );
  Memory_198 rotation45deg_33 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_33_clock),
    .io_address(rotation45deg_33_io_address)
  );
  Memory_198 rotation45deg_34 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_34_clock),
    .io_address(rotation45deg_34_io_address)
  );
  Memory_198 rotation45deg_35 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_35_clock),
    .io_address(rotation45deg_35_io_address)
  );
  Memory_198 rotation45deg_36 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_36_clock),
    .io_address(rotation45deg_36_io_address)
  );
  Memory_198 rotation45deg_37 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_37_clock),
    .io_address(rotation45deg_37_io_address)
  );
  Memory_198 rotation45deg_38 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_38_clock),
    .io_address(rotation45deg_38_io_address)
  );
  Memory_198 rotation45deg_39 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_39_clock),
    .io_address(rotation45deg_39_io_address)
  );
  Memory_198 rotation45deg_40 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_40_clock),
    .io_address(rotation45deg_40_io_address)
  );
  Memory_198 rotation45deg_41 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_41_clock),
    .io_address(rotation45deg_41_io_address)
  );
  Memory_198 rotation45deg_42 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_42_clock),
    .io_address(rotation45deg_42_io_address)
  );
  Memory_198 rotation45deg_43 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_43_clock),
    .io_address(rotation45deg_43_io_address)
  );
  Memory_198 rotation45deg_44 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_44_clock),
    .io_address(rotation45deg_44_io_address)
  );
  Memory_198 rotation45deg_45 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_45_clock),
    .io_address(rotation45deg_45_io_address)
  );
  Memory_198 rotation45deg_46 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_46_clock),
    .io_address(rotation45deg_46_io_address)
  );
  Memory_198 rotation45deg_47 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_47_clock),
    .io_address(rotation45deg_47_io_address)
  );
  Memory_198 rotation45deg_48 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_48_clock),
    .io_address(rotation45deg_48_io_address)
  );
  Memory_198 rotation45deg_49 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_49_clock),
    .io_address(rotation45deg_49_io_address)
  );
  Memory_198 rotation45deg_50 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_50_clock),
    .io_address(rotation45deg_50_io_address)
  );
  Memory_198 rotation45deg_51 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_51_clock),
    .io_address(rotation45deg_51_io_address)
  );
  Memory_198 rotation45deg_52 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_52_clock),
    .io_address(rotation45deg_52_io_address)
  );
  Memory_198 rotation45deg_53 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_53_clock),
    .io_address(rotation45deg_53_io_address)
  );
  Memory_198 rotation45deg_54 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_54_clock),
    .io_address(rotation45deg_54_io_address)
  );
  Memory_198 rotation45deg_55 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_55_clock),
    .io_address(rotation45deg_55_io_address)
  );
  Memory_198 rotation45deg_56 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_56_clock),
    .io_address(rotation45deg_56_io_address)
  );
  Memory_198 rotation45deg_57 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_57_clock),
    .io_address(rotation45deg_57_io_address)
  );
  Memory_198 rotation45deg_58 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_58_clock),
    .io_address(rotation45deg_58_io_address)
  );
  Memory_198 rotation45deg_59 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_59_clock),
    .io_address(rotation45deg_59_io_address)
  );
  Memory_198 rotation45deg_60 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_60_clock),
    .io_address(rotation45deg_60_io_address)
  );
  Memory_198 rotation45deg_61 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_61_clock),
    .io_address(rotation45deg_61_io_address)
  );
  Memory_198 rotation45deg_62 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_62_clock),
    .io_address(rotation45deg_62_io_address)
  );
  Memory_198 rotation45deg_63 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_63_clock),
    .io_address(rotation45deg_63_io_address)
  );
  Memory_198 rotation45deg_64 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_64_clock),
    .io_address(rotation45deg_64_io_address)
  );
  Memory_198 rotation45deg_65 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_65_clock),
    .io_address(rotation45deg_65_io_address)
  );
  Memory_198 rotation45deg_66 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_66_clock),
    .io_address(rotation45deg_66_io_address)
  );
  Memory_198 rotation45deg_67 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_67_clock),
    .io_address(rotation45deg_67_io_address)
  );
  Memory_198 rotation45deg_68 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_68_clock),
    .io_address(rotation45deg_68_io_address)
  );
  Memory_198 rotation45deg_69 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_69_clock),
    .io_address(rotation45deg_69_io_address)
  );
  Memory_198 rotation45deg_70 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_70_clock),
    .io_address(rotation45deg_70_io_address)
  );
  Memory_198 rotation45deg_71 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_71_clock),
    .io_address(rotation45deg_71_io_address)
  );
  Memory_198 rotation45deg_72 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_72_clock),
    .io_address(rotation45deg_72_io_address)
  );
  Memory_198 rotation45deg_73 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_73_clock),
    .io_address(rotation45deg_73_io_address)
  );
  Memory_198 rotation45deg_74 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_74_clock),
    .io_address(rotation45deg_74_io_address)
  );
  Memory_198 rotation45deg_75 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_75_clock),
    .io_address(rotation45deg_75_io_address)
  );
  Memory_198 rotation45deg_76 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_76_clock),
    .io_address(rotation45deg_76_io_address)
  );
  Memory_198 rotation45deg_77 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_77_clock),
    .io_address(rotation45deg_77_io_address)
  );
  Memory_198 rotation45deg_78 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_78_clock),
    .io_address(rotation45deg_78_io_address)
  );
  Memory_198 rotation45deg_79 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_79_clock),
    .io_address(rotation45deg_79_io_address)
  );
  Memory_198 rotation45deg_80 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_80_clock),
    .io_address(rotation45deg_80_io_address)
  );
  Memory_198 rotation45deg_81 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_81_clock),
    .io_address(rotation45deg_81_io_address)
  );
  Memory_198 rotation45deg_82 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_82_clock),
    .io_address(rotation45deg_82_io_address)
  );
  Memory_198 rotation45deg_83 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_83_clock),
    .io_address(rotation45deg_83_io_address)
  );
  Memory_198 rotation45deg_84 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_84_clock),
    .io_address(rotation45deg_84_io_address)
  );
  Memory_198 rotation45deg_85 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_85_clock),
    .io_address(rotation45deg_85_io_address)
  );
  Memory_198 rotation45deg_86 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_86_clock),
    .io_address(rotation45deg_86_io_address)
  );
  Memory_198 rotation45deg_87 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_87_clock),
    .io_address(rotation45deg_87_io_address)
  );
  Memory_198 rotation45deg_88 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_88_clock),
    .io_address(rotation45deg_88_io_address)
  );
  Memory_198 rotation45deg_89 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_89_clock),
    .io_address(rotation45deg_89_io_address)
  );
  Memory_198 rotation45deg_90 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_90_clock),
    .io_address(rotation45deg_90_io_address)
  );
  Memory_198 rotation45deg_91 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_91_clock),
    .io_address(rotation45deg_91_io_address)
  );
  Memory_198 rotation45deg_92 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_92_clock),
    .io_address(rotation45deg_92_io_address)
  );
  Memory_198 rotation45deg_93 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_93_clock),
    .io_address(rotation45deg_93_io_address)
  );
  Memory_198 rotation45deg_94 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_94_clock),
    .io_address(rotation45deg_94_io_address)
  );
  Memory_198 rotation45deg_95 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_95_clock),
    .io_address(rotation45deg_95_io_address)
  );
  Memory_198 rotation45deg_96 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_96_clock),
    .io_address(rotation45deg_96_io_address)
  );
  Memory_198 rotation45deg_97 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_97_clock),
    .io_address(rotation45deg_97_io_address)
  );
  Memory_198 rotation45deg_98 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_98_clock),
    .io_address(rotation45deg_98_io_address)
  );
  Memory_198 rotation45deg_99 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_99_clock),
    .io_address(rotation45deg_99_io_address)
  );
  Memory_198 rotation45deg_100 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_100_clock),
    .io_address(rotation45deg_100_io_address)
  );
  Memory_198 rotation45deg_101 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_101_clock),
    .io_address(rotation45deg_101_io_address)
  );
  Memory_198 rotation45deg_102 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_102_clock),
    .io_address(rotation45deg_102_io_address)
  );
  Memory_198 rotation45deg_103 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_103_clock),
    .io_address(rotation45deg_103_io_address)
  );
  Memory_198 rotation45deg_104 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_104_clock),
    .io_address(rotation45deg_104_io_address)
  );
  Memory_198 rotation45deg_105 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_105_clock),
    .io_address(rotation45deg_105_io_address)
  );
  Memory_198 rotation45deg_106 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_106_clock),
    .io_address(rotation45deg_106_io_address)
  );
  Memory_198 rotation45deg_107 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_107_clock),
    .io_address(rotation45deg_107_io_address)
  );
  Memory_198 rotation45deg_108 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_108_clock),
    .io_address(rotation45deg_108_io_address)
  );
  Memory_198 rotation45deg_109 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_109_clock),
    .io_address(rotation45deg_109_io_address)
  );
  Memory_198 rotation45deg_110 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_110_clock),
    .io_address(rotation45deg_110_io_address)
  );
  Memory_198 rotation45deg_111 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_111_clock),
    .io_address(rotation45deg_111_io_address)
  );
  Memory_198 rotation45deg_112 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_112_clock),
    .io_address(rotation45deg_112_io_address)
  );
  Memory_198 rotation45deg_113 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_113_clock),
    .io_address(rotation45deg_113_io_address)
  );
  Memory_198 rotation45deg_114 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_114_clock),
    .io_address(rotation45deg_114_io_address)
  );
  Memory_198 rotation45deg_115 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_115_clock),
    .io_address(rotation45deg_115_io_address)
  );
  Memory_198 rotation45deg_116 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_116_clock),
    .io_address(rotation45deg_116_io_address)
  );
  Memory_198 rotation45deg_117 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_117_clock),
    .io_address(rotation45deg_117_io_address)
  );
  Memory_198 rotation45deg_118 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_118_clock),
    .io_address(rotation45deg_118_io_address)
  );
  Memory_198 rotation45deg_119 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_119_clock),
    .io_address(rotation45deg_119_io_address)
  );
  Memory_198 rotation45deg_120 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_120_clock),
    .io_address(rotation45deg_120_io_address)
  );
  Memory_198 rotation45deg_121 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_121_clock),
    .io_address(rotation45deg_121_io_address)
  );
  Memory_198 rotation45deg_122 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_122_clock),
    .io_address(rotation45deg_122_io_address)
  );
  Memory_198 rotation45deg_123 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_123_clock),
    .io_address(rotation45deg_123_io_address)
  );
  Memory_198 rotation45deg_124 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_124_clock),
    .io_address(rotation45deg_124_io_address)
  );
  Memory_198 rotation45deg_125 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_125_clock),
    .io_address(rotation45deg_125_io_address)
  );
  Memory_198 rotation45deg_126 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_126_clock),
    .io_address(rotation45deg_126_io_address)
  );
  Memory_198 rotation45deg_127 ( // @[GraphicEngineVGA.scala 325:30]
    .clock(rotation45deg_127_clock),
    .io_address(rotation45deg_127_io_address)
  );
  SpriteBlender spriteBlender ( // @[GraphicEngineVGA.scala 333:29]
    .clock(spriteBlender_clock),
    .io_pixelColorBack(spriteBlender_io_pixelColorBack),
    .io_spriteVisibleReg_0(spriteBlender_io_spriteVisibleReg_0),
    .io_spriteVisibleReg_1(spriteBlender_io_spriteVisibleReg_1),
    .io_spriteVisibleReg_2(spriteBlender_io_spriteVisibleReg_2),
    .io_spriteVisibleReg_3(spriteBlender_io_spriteVisibleReg_3),
    .io_spriteVisibleReg_4(spriteBlender_io_spriteVisibleReg_4),
    .io_spriteVisibleReg_5(spriteBlender_io_spriteVisibleReg_5),
    .io_spriteVisibleReg_6(spriteBlender_io_spriteVisibleReg_6),
    .io_spriteVisibleReg_7(spriteBlender_io_spriteVisibleReg_7),
    .io_spriteVisibleReg_8(spriteBlender_io_spriteVisibleReg_8),
    .io_spriteVisibleReg_9(spriteBlender_io_spriteVisibleReg_9),
    .io_spriteVisibleReg_10(spriteBlender_io_spriteVisibleReg_10),
    .io_spriteVisibleReg_11(spriteBlender_io_spriteVisibleReg_11),
    .io_spriteVisibleReg_12(spriteBlender_io_spriteVisibleReg_12),
    .io_spriteVisibleReg_13(spriteBlender_io_spriteVisibleReg_13),
    .io_spriteVisibleReg_14(spriteBlender_io_spriteVisibleReg_14),
    .io_spriteVisibleReg_15(spriteBlender_io_spriteVisibleReg_15),
    .io_spriteVisibleReg_16(spriteBlender_io_spriteVisibleReg_16),
    .io_spriteVisibleReg_17(spriteBlender_io_spriteVisibleReg_17),
    .io_spriteVisibleReg_18(spriteBlender_io_spriteVisibleReg_18),
    .io_spriteVisibleReg_19(spriteBlender_io_spriteVisibleReg_19),
    .io_spriteVisibleReg_20(spriteBlender_io_spriteVisibleReg_20),
    .io_spriteVisibleReg_21(spriteBlender_io_spriteVisibleReg_21),
    .io_spriteVisibleReg_22(spriteBlender_io_spriteVisibleReg_22),
    .io_spriteVisibleReg_23(spriteBlender_io_spriteVisibleReg_23),
    .io_spriteVisibleReg_24(spriteBlender_io_spriteVisibleReg_24),
    .io_spriteVisibleReg_25(spriteBlender_io_spriteVisibleReg_25),
    .io_spriteVisibleReg_26(spriteBlender_io_spriteVisibleReg_26),
    .io_spriteVisibleReg_27(spriteBlender_io_spriteVisibleReg_27),
    .io_spriteVisibleReg_28(spriteBlender_io_spriteVisibleReg_28),
    .io_spriteVisibleReg_29(spriteBlender_io_spriteVisibleReg_29),
    .io_spriteVisibleReg_30(spriteBlender_io_spriteVisibleReg_30),
    .io_spriteVisibleReg_31(spriteBlender_io_spriteVisibleReg_31),
    .io_spriteVisibleReg_32(spriteBlender_io_spriteVisibleReg_32),
    .io_spriteVisibleReg_33(spriteBlender_io_spriteVisibleReg_33),
    .io_spriteVisibleReg_41(spriteBlender_io_spriteVisibleReg_41),
    .io_spriteVisibleReg_42(spriteBlender_io_spriteVisibleReg_42),
    .io_spriteVisibleReg_43(spriteBlender_io_spriteVisibleReg_43),
    .io_spriteVisibleReg_44(spriteBlender_io_spriteVisibleReg_44),
    .io_spriteVisibleReg_45(spriteBlender_io_spriteVisibleReg_45),
    .io_spriteVisibleReg_46(spriteBlender_io_spriteVisibleReg_46),
    .io_spriteVisibleReg_47(spriteBlender_io_spriteVisibleReg_47),
    .io_spriteVisibleReg_48(spriteBlender_io_spriteVisibleReg_48),
    .io_spriteVisibleReg_49(spriteBlender_io_spriteVisibleReg_49),
    .io_spriteVisibleReg_50(spriteBlender_io_spriteVisibleReg_50),
    .io_spriteVisibleReg_51(spriteBlender_io_spriteVisibleReg_51),
    .io_spriteVisibleReg_55(spriteBlender_io_spriteVisibleReg_55),
    .io_spriteVisibleReg_56(spriteBlender_io_spriteVisibleReg_56),
    .io_spriteVisibleReg_57(spriteBlender_io_spriteVisibleReg_57),
    .io_spriteVisibleReg_61(spriteBlender_io_spriteVisibleReg_61),
    .io_spriteVisibleReg_62(spriteBlender_io_spriteVisibleReg_62),
    .io_spriteVisibleReg_63(spriteBlender_io_spriteVisibleReg_63),
    .io_spriteVisibleReg_64(spriteBlender_io_spriteVisibleReg_64),
    .io_spriteVisibleReg_65(spriteBlender_io_spriteVisibleReg_65),
    .io_spriteVisibleReg_66(spriteBlender_io_spriteVisibleReg_66),
    .io_spriteVisibleReg_70(spriteBlender_io_spriteVisibleReg_70),
    .io_spriteVisibleReg_71(spriteBlender_io_spriteVisibleReg_71),
    .io_spriteVisibleReg_72(spriteBlender_io_spriteVisibleReg_72),
    .io_inSprite_0(spriteBlender_io_inSprite_0),
    .io_inSprite_1(spriteBlender_io_inSprite_1),
    .io_inSprite_2(spriteBlender_io_inSprite_2),
    .io_inSprite_3(spriteBlender_io_inSprite_3),
    .io_inSprite_4(spriteBlender_io_inSprite_4),
    .io_inSprite_5(spriteBlender_io_inSprite_5),
    .io_inSprite_6(spriteBlender_io_inSprite_6),
    .io_inSprite_7(spriteBlender_io_inSprite_7),
    .io_inSprite_8(spriteBlender_io_inSprite_8),
    .io_inSprite_9(spriteBlender_io_inSprite_9),
    .io_inSprite_10(spriteBlender_io_inSprite_10),
    .io_inSprite_11(spriteBlender_io_inSprite_11),
    .io_inSprite_12(spriteBlender_io_inSprite_12),
    .io_inSprite_13(spriteBlender_io_inSprite_13),
    .io_inSprite_14(spriteBlender_io_inSprite_14),
    .io_inSprite_15(spriteBlender_io_inSprite_15),
    .io_inSprite_16(spriteBlender_io_inSprite_16),
    .io_inSprite_17(spriteBlender_io_inSprite_17),
    .io_inSprite_18(spriteBlender_io_inSprite_18),
    .io_inSprite_19(spriteBlender_io_inSprite_19),
    .io_inSprite_20(spriteBlender_io_inSprite_20),
    .io_inSprite_21(spriteBlender_io_inSprite_21),
    .io_inSprite_22(spriteBlender_io_inSprite_22),
    .io_inSprite_23(spriteBlender_io_inSprite_23),
    .io_inSprite_24(spriteBlender_io_inSprite_24),
    .io_inSprite_25(spriteBlender_io_inSprite_25),
    .io_inSprite_26(spriteBlender_io_inSprite_26),
    .io_inSprite_27(spriteBlender_io_inSprite_27),
    .io_inSprite_28(spriteBlender_io_inSprite_28),
    .io_inSprite_29(spriteBlender_io_inSprite_29),
    .io_inSprite_30(spriteBlender_io_inSprite_30),
    .io_inSprite_31(spriteBlender_io_inSprite_31),
    .io_inSprite_32(spriteBlender_io_inSprite_32),
    .io_inSprite_33(spriteBlender_io_inSprite_33),
    .io_inSprite_34(spriteBlender_io_inSprite_34),
    .io_inSprite_35(spriteBlender_io_inSprite_35),
    .io_inSprite_36(spriteBlender_io_inSprite_36),
    .io_inSprite_37(spriteBlender_io_inSprite_37),
    .io_inSprite_38(spriteBlender_io_inSprite_38),
    .io_inSprite_39(spriteBlender_io_inSprite_39),
    .io_inSprite_40(spriteBlender_io_inSprite_40),
    .io_inSprite_41(spriteBlender_io_inSprite_41),
    .io_inSprite_42(spriteBlender_io_inSprite_42),
    .io_inSprite_43(spriteBlender_io_inSprite_43),
    .io_inSprite_44(spriteBlender_io_inSprite_44),
    .io_inSprite_45(spriteBlender_io_inSprite_45),
    .io_inSprite_46(spriteBlender_io_inSprite_46),
    .io_inSprite_47(spriteBlender_io_inSprite_47),
    .io_inSprite_48(spriteBlender_io_inSprite_48),
    .io_inSprite_49(spriteBlender_io_inSprite_49),
    .io_inSprite_50(spriteBlender_io_inSprite_50),
    .io_inSprite_51(spriteBlender_io_inSprite_51),
    .io_inSprite_52(spriteBlender_io_inSprite_52),
    .io_inSprite_53(spriteBlender_io_inSprite_53),
    .io_inSprite_54(spriteBlender_io_inSprite_54),
    .io_inSprite_55(spriteBlender_io_inSprite_55),
    .io_inSprite_56(spriteBlender_io_inSprite_56),
    .io_inSprite_57(spriteBlender_io_inSprite_57),
    .io_inSprite_58(spriteBlender_io_inSprite_58),
    .io_inSprite_59(spriteBlender_io_inSprite_59),
    .io_inSprite_60(spriteBlender_io_inSprite_60),
    .io_inSprite_61(spriteBlender_io_inSprite_61),
    .io_inSprite_62(spriteBlender_io_inSprite_62),
    .io_inSprite_63(spriteBlender_io_inSprite_63),
    .io_inSprite_64(spriteBlender_io_inSprite_64),
    .io_inSprite_65(spriteBlender_io_inSprite_65),
    .io_inSprite_66(spriteBlender_io_inSprite_66),
    .io_inSprite_67(spriteBlender_io_inSprite_67),
    .io_inSprite_68(spriteBlender_io_inSprite_68),
    .io_inSprite_69(spriteBlender_io_inSprite_69),
    .io_inSprite_70(spriteBlender_io_inSprite_70),
    .io_inSprite_71(spriteBlender_io_inSprite_71),
    .io_inSprite_72(spriteBlender_io_inSprite_72),
    .io_inSprite_73(spriteBlender_io_inSprite_73),
    .io_inSprite_74(spriteBlender_io_inSprite_74),
    .io_inSprite_75(spriteBlender_io_inSprite_75),
    .io_inSprite_76(spriteBlender_io_inSprite_76),
    .io_inSprite_77(spriteBlender_io_inSprite_77),
    .io_inSprite_78(spriteBlender_io_inSprite_78),
    .io_inSprite_79(spriteBlender_io_inSprite_79),
    .io_inSprite_80(spriteBlender_io_inSprite_80),
    .io_inSprite_81(spriteBlender_io_inSprite_81),
    .io_inSprite_82(spriteBlender_io_inSprite_82),
    .io_inSprite_83(spriteBlender_io_inSprite_83),
    .io_inSprite_84(spriteBlender_io_inSprite_84),
    .io_inSprite_85(spriteBlender_io_inSprite_85),
    .io_inSprite_86(spriteBlender_io_inSprite_86),
    .io_inSprite_87(spriteBlender_io_inSprite_87),
    .io_inSprite_88(spriteBlender_io_inSprite_88),
    .io_inSprite_89(spriteBlender_io_inSprite_89),
    .io_inSprite_90(spriteBlender_io_inSprite_90),
    .io_inSprite_91(spriteBlender_io_inSprite_91),
    .io_inSprite_92(spriteBlender_io_inSprite_92),
    .io_inSprite_93(spriteBlender_io_inSprite_93),
    .io_inSprite_94(spriteBlender_io_inSprite_94),
    .io_inSprite_95(spriteBlender_io_inSprite_95),
    .io_inSprite_96(spriteBlender_io_inSprite_96),
    .io_inSprite_97(spriteBlender_io_inSprite_97),
    .io_inSprite_98(spriteBlender_io_inSprite_98),
    .io_inSprite_99(spriteBlender_io_inSprite_99),
    .io_inSprite_100(spriteBlender_io_inSprite_100),
    .io_inSprite_101(spriteBlender_io_inSprite_101),
    .io_inSprite_102(spriteBlender_io_inSprite_102),
    .io_inSprite_103(spriteBlender_io_inSprite_103),
    .io_inSprite_104(spriteBlender_io_inSprite_104),
    .io_inSprite_105(spriteBlender_io_inSprite_105),
    .io_inSprite_106(spriteBlender_io_inSprite_106),
    .io_inSprite_107(spriteBlender_io_inSprite_107),
    .io_inSprite_108(spriteBlender_io_inSprite_108),
    .io_inSprite_109(spriteBlender_io_inSprite_109),
    .io_inSprite_110(spriteBlender_io_inSprite_110),
    .io_inSprite_111(spriteBlender_io_inSprite_111),
    .io_inSprite_112(spriteBlender_io_inSprite_112),
    .io_inSprite_113(spriteBlender_io_inSprite_113),
    .io_inSprite_114(spriteBlender_io_inSprite_114),
    .io_inSprite_115(spriteBlender_io_inSprite_115),
    .io_inSprite_116(spriteBlender_io_inSprite_116),
    .io_inSprite_117(spriteBlender_io_inSprite_117),
    .io_inSprite_118(spriteBlender_io_inSprite_118),
    .io_inSprite_119(spriteBlender_io_inSprite_119),
    .io_inSprite_120(spriteBlender_io_inSprite_120),
    .io_inSprite_121(spriteBlender_io_inSprite_121),
    .io_inSprite_122(spriteBlender_io_inSprite_122),
    .io_inSprite_123(spriteBlender_io_inSprite_123),
    .io_inSprite_124(spriteBlender_io_inSprite_124),
    .io_inSprite_125(spriteBlender_io_inSprite_125),
    .io_inSprite_126(spriteBlender_io_inSprite_126),
    .io_inSprite_127(spriteBlender_io_inSprite_127),
    .io_datareader_0(spriteBlender_io_datareader_0),
    .io_datareader_1(spriteBlender_io_datareader_1),
    .io_datareader_2(spriteBlender_io_datareader_2),
    .io_datareader_3(spriteBlender_io_datareader_3),
    .io_datareader_4(spriteBlender_io_datareader_4),
    .io_datareader_5(spriteBlender_io_datareader_5),
    .io_datareader_6(spriteBlender_io_datareader_6),
    .io_datareader_7(spriteBlender_io_datareader_7),
    .io_datareader_8(spriteBlender_io_datareader_8),
    .io_datareader_9(spriteBlender_io_datareader_9),
    .io_datareader_10(spriteBlender_io_datareader_10),
    .io_datareader_11(spriteBlender_io_datareader_11),
    .io_datareader_12(spriteBlender_io_datareader_12),
    .io_datareader_13(spriteBlender_io_datareader_13),
    .io_datareader_14(spriteBlender_io_datareader_14),
    .io_datareader_15(spriteBlender_io_datareader_15),
    .io_datareader_16(spriteBlender_io_datareader_16),
    .io_datareader_17(spriteBlender_io_datareader_17),
    .io_datareader_18(spriteBlender_io_datareader_18),
    .io_datareader_19(spriteBlender_io_datareader_19),
    .io_datareader_20(spriteBlender_io_datareader_20),
    .io_datareader_21(spriteBlender_io_datareader_21),
    .io_datareader_22(spriteBlender_io_datareader_22),
    .io_datareader_23(spriteBlender_io_datareader_23),
    .io_datareader_24(spriteBlender_io_datareader_24),
    .io_datareader_25(spriteBlender_io_datareader_25),
    .io_datareader_26(spriteBlender_io_datareader_26),
    .io_datareader_27(spriteBlender_io_datareader_27),
    .io_datareader_28(spriteBlender_io_datareader_28),
    .io_datareader_29(spriteBlender_io_datareader_29),
    .io_datareader_30(spriteBlender_io_datareader_30),
    .io_datareader_31(spriteBlender_io_datareader_31),
    .io_datareader_32(spriteBlender_io_datareader_32),
    .io_datareader_33(spriteBlender_io_datareader_33),
    .io_datareader_34(spriteBlender_io_datareader_34),
    .io_datareader_35(spriteBlender_io_datareader_35),
    .io_datareader_36(spriteBlender_io_datareader_36),
    .io_datareader_37(spriteBlender_io_datareader_37),
    .io_datareader_38(spriteBlender_io_datareader_38),
    .io_datareader_39(spriteBlender_io_datareader_39),
    .io_datareader_40(spriteBlender_io_datareader_40),
    .io_datareader_41(spriteBlender_io_datareader_41),
    .io_datareader_42(spriteBlender_io_datareader_42),
    .io_datareader_43(spriteBlender_io_datareader_43),
    .io_datareader_44(spriteBlender_io_datareader_44),
    .io_datareader_45(spriteBlender_io_datareader_45),
    .io_datareader_46(spriteBlender_io_datareader_46),
    .io_datareader_47(spriteBlender_io_datareader_47),
    .io_datareader_48(spriteBlender_io_datareader_48),
    .io_datareader_49(spriteBlender_io_datareader_49),
    .io_datareader_50(spriteBlender_io_datareader_50),
    .io_datareader_51(spriteBlender_io_datareader_51),
    .io_datareader_52(spriteBlender_io_datareader_52),
    .io_datareader_53(spriteBlender_io_datareader_53),
    .io_datareader_54(spriteBlender_io_datareader_54),
    .io_datareader_55(spriteBlender_io_datareader_55),
    .io_datareader_56(spriteBlender_io_datareader_56),
    .io_datareader_57(spriteBlender_io_datareader_57),
    .io_datareader_58(spriteBlender_io_datareader_58),
    .io_datareader_59(spriteBlender_io_datareader_59),
    .io_datareader_60(spriteBlender_io_datareader_60),
    .io_datareader_61(spriteBlender_io_datareader_61),
    .io_datareader_62(spriteBlender_io_datareader_62),
    .io_datareader_63(spriteBlender_io_datareader_63),
    .io_datareader_64(spriteBlender_io_datareader_64),
    .io_datareader_65(spriteBlender_io_datareader_65),
    .io_datareader_66(spriteBlender_io_datareader_66),
    .io_datareader_67(spriteBlender_io_datareader_67),
    .io_datareader_68(spriteBlender_io_datareader_68),
    .io_datareader_69(spriteBlender_io_datareader_69),
    .io_datareader_70(spriteBlender_io_datareader_70),
    .io_datareader_71(spriteBlender_io_datareader_71),
    .io_datareader_72(spriteBlender_io_datareader_72),
    .io_datareader_73(spriteBlender_io_datareader_73),
    .io_datareader_74(spriteBlender_io_datareader_74),
    .io_datareader_75(spriteBlender_io_datareader_75),
    .io_datareader_76(spriteBlender_io_datareader_76),
    .io_datareader_77(spriteBlender_io_datareader_77),
    .io_datareader_78(spriteBlender_io_datareader_78),
    .io_datareader_79(spriteBlender_io_datareader_79),
    .io_datareader_80(spriteBlender_io_datareader_80),
    .io_datareader_81(spriteBlender_io_datareader_81),
    .io_datareader_82(spriteBlender_io_datareader_82),
    .io_datareader_83(spriteBlender_io_datareader_83),
    .io_datareader_84(spriteBlender_io_datareader_84),
    .io_datareader_85(spriteBlender_io_datareader_85),
    .io_datareader_86(spriteBlender_io_datareader_86),
    .io_datareader_87(spriteBlender_io_datareader_87),
    .io_datareader_88(spriteBlender_io_datareader_88),
    .io_datareader_89(spriteBlender_io_datareader_89),
    .io_datareader_90(spriteBlender_io_datareader_90),
    .io_datareader_91(spriteBlender_io_datareader_91),
    .io_datareader_92(spriteBlender_io_datareader_92),
    .io_datareader_93(spriteBlender_io_datareader_93),
    .io_datareader_94(spriteBlender_io_datareader_94),
    .io_datareader_95(spriteBlender_io_datareader_95),
    .io_datareader_96(spriteBlender_io_datareader_96),
    .io_datareader_97(spriteBlender_io_datareader_97),
    .io_datareader_98(spriteBlender_io_datareader_98),
    .io_datareader_99(spriteBlender_io_datareader_99),
    .io_datareader_100(spriteBlender_io_datareader_100),
    .io_datareader_101(spriteBlender_io_datareader_101),
    .io_datareader_102(spriteBlender_io_datareader_102),
    .io_datareader_103(spriteBlender_io_datareader_103),
    .io_datareader_104(spriteBlender_io_datareader_104),
    .io_datareader_105(spriteBlender_io_datareader_105),
    .io_datareader_106(spriteBlender_io_datareader_106),
    .io_datareader_107(spriteBlender_io_datareader_107),
    .io_datareader_108(spriteBlender_io_datareader_108),
    .io_datareader_109(spriteBlender_io_datareader_109),
    .io_datareader_110(spriteBlender_io_datareader_110),
    .io_datareader_111(spriteBlender_io_datareader_111),
    .io_datareader_112(spriteBlender_io_datareader_112),
    .io_datareader_113(spriteBlender_io_datareader_113),
    .io_datareader_114(spriteBlender_io_datareader_114),
    .io_datareader_115(spriteBlender_io_datareader_115),
    .io_datareader_116(spriteBlender_io_datareader_116),
    .io_datareader_117(spriteBlender_io_datareader_117),
    .io_datareader_118(spriteBlender_io_datareader_118),
    .io_datareader_119(spriteBlender_io_datareader_119),
    .io_datareader_120(spriteBlender_io_datareader_120),
    .io_datareader_121(spriteBlender_io_datareader_121),
    .io_datareader_122(spriteBlender_io_datareader_122),
    .io_datareader_123(spriteBlender_io_datareader_123),
    .io_datareader_124(spriteBlender_io_datareader_124),
    .io_datareader_125(spriteBlender_io_datareader_125),
    .io_datareader_126(spriteBlender_io_datareader_126),
    .io_datareader_127(spriteBlender_io_datareader_127),
    .io_vgaRed(spriteBlender_io_vgaRed),
    .io_vgaGreen(spriteBlender_io_vgaGreen),
    .io_vgaBlue(spriteBlender_io_vgaBlue)
  );
  assign io_newFrame = run & _GEN_8; // @[GraphicEngineVGA.scala 78:15 GraphicEngineVGA.scala 88:23]
  assign io_missingFrameError = missingFrameErrorReg; // @[GraphicEngineVGA.scala 149:24]
  assign io_backBufferWriteError = backBufferWriteErrorReg; // @[GraphicEngineVGA.scala 150:27]
  assign io_viewBoxOutOfRangeError = viewBoxOutOfRangeErrorReg; // @[GraphicEngineVGA.scala 151:29]
  assign io_vgaRed = _T_15660_0 ? spriteBlender_io_vgaRed : 4'h0; // @[GraphicEngineVGA.scala 412:13 GraphicEngineVGA.scala 416:13]
  assign io_vgaBlue = _T_15664_0 ? spriteBlender_io_vgaBlue : 4'h0; // @[GraphicEngineVGA.scala 413:14 GraphicEngineVGA.scala 418:13]
  assign io_vgaGreen = _T_15662_0 ? spriteBlender_io_vgaGreen : 4'h0; // @[GraphicEngineVGA.scala 414:15 GraphicEngineVGA.scala 417:14]
  assign io_Hsync = _T_14_0; // @[GraphicEngineVGA.scala 102:12]
  assign io_Vsync = _T_16_0; // @[GraphicEngineVGA.scala 103:12]
  assign backTileMemories_0_0_clock = clock;
  assign backTileMemories_0_0_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_1_clock = clock;
  assign backTileMemories_0_1_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_2_clock = clock;
  assign backTileMemories_0_2_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_3_clock = clock;
  assign backTileMemories_0_3_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_4_clock = clock;
  assign backTileMemories_0_4_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_5_clock = clock;
  assign backTileMemories_0_5_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_6_clock = clock;
  assign backTileMemories_0_6_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_7_clock = clock;
  assign backTileMemories_0_7_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_8_clock = clock;
  assign backTileMemories_0_8_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_9_clock = clock;
  assign backTileMemories_0_9_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_10_clock = clock;
  assign backTileMemories_0_10_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_11_clock = clock;
  assign backTileMemories_0_11_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_12_clock = clock;
  assign backTileMemories_0_12_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_13_clock = clock;
  assign backTileMemories_0_13_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_14_clock = clock;
  assign backTileMemories_0_14_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_15_clock = clock;
  assign backTileMemories_0_15_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_16_clock = clock;
  assign backTileMemories_0_16_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_17_clock = clock;
  assign backTileMemories_0_17_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_18_clock = clock;
  assign backTileMemories_0_18_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_19_clock = clock;
  assign backTileMemories_0_19_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_20_clock = clock;
  assign backTileMemories_0_20_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_21_clock = clock;
  assign backTileMemories_0_21_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_22_clock = clock;
  assign backTileMemories_0_22_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_23_clock = clock;
  assign backTileMemories_0_23_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_24_clock = clock;
  assign backTileMemories_0_24_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_25_clock = clock;
  assign backTileMemories_0_25_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_26_clock = clock;
  assign backTileMemories_0_26_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_27_clock = clock;
  assign backTileMemories_0_27_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_28_clock = clock;
  assign backTileMemories_0_28_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_29_clock = clock;
  assign backTileMemories_0_29_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_30_clock = clock;
  assign backTileMemories_0_30_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_0_31_clock = clock;
  assign backTileMemories_0_31_io_address = _T_52[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_0_clock = clock;
  assign backTileMemories_1_0_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_1_clock = clock;
  assign backTileMemories_1_1_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_2_clock = clock;
  assign backTileMemories_1_2_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_3_clock = clock;
  assign backTileMemories_1_3_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_4_clock = clock;
  assign backTileMemories_1_4_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_5_clock = clock;
  assign backTileMemories_1_5_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_6_clock = clock;
  assign backTileMemories_1_6_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_7_clock = clock;
  assign backTileMemories_1_7_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_8_clock = clock;
  assign backTileMemories_1_8_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_9_clock = clock;
  assign backTileMemories_1_9_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_10_clock = clock;
  assign backTileMemories_1_10_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_11_clock = clock;
  assign backTileMemories_1_11_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_12_clock = clock;
  assign backTileMemories_1_12_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_13_clock = clock;
  assign backTileMemories_1_13_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_14_clock = clock;
  assign backTileMemories_1_14_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_15_clock = clock;
  assign backTileMemories_1_15_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_16_clock = clock;
  assign backTileMemories_1_16_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_17_clock = clock;
  assign backTileMemories_1_17_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_18_clock = clock;
  assign backTileMemories_1_18_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_19_clock = clock;
  assign backTileMemories_1_19_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_20_clock = clock;
  assign backTileMemories_1_20_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_21_clock = clock;
  assign backTileMemories_1_21_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_22_clock = clock;
  assign backTileMemories_1_22_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_23_clock = clock;
  assign backTileMemories_1_23_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_24_clock = clock;
  assign backTileMemories_1_24_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_25_clock = clock;
  assign backTileMemories_1_25_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_26_clock = clock;
  assign backTileMemories_1_26_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_27_clock = clock;
  assign backTileMemories_1_27_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_28_clock = clock;
  assign backTileMemories_1_28_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_29_clock = clock;
  assign backTileMemories_1_29_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_30_clock = clock;
  assign backTileMemories_1_30_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backTileMemories_1_31_clock = clock;
  assign backTileMemories_1_31_io_address = _T_212[9:0]; // @[GraphicEngineVGA.scala 220:39]
  assign backBufferMemories_0_clock = clock;
  assign backBufferMemories_0_io_address = _T_394[10:0]; // @[GraphicEngineVGA.scala 292:36]
  assign backBufferMemories_0_io_writeEnable = copyEnabledReg; // @[GraphicEngineVGA.scala 294:40]
  assign backBufferMemories_0_io_dataWrite = backBufferShadowMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 295:38]
  assign backBufferMemories_1_clock = clock;
  assign backBufferMemories_1_io_address = _T_414[10:0]; // @[GraphicEngineVGA.scala 292:36]
  assign backBufferMemories_1_io_writeEnable = copyEnabledReg; // @[GraphicEngineVGA.scala 294:40]
  assign backBufferMemories_1_io_dataWrite = backBufferShadowMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 295:38]
  assign backBufferShadowMemories_0_clock = clock;
  assign backBufferShadowMemories_0_io_address = restoreEnabled ? _T_377 : _T_380; // @[GraphicEngineVGA.scala 287:42]
  assign backBufferShadowMemories_0_io_writeEnable = restoreEnabled ? _T_382 : _T_384; // @[GraphicEngineVGA.scala 289:46]
  assign backBufferShadowMemories_0_io_dataWrite = restoreEnabled ? backBufferRestoreMemories_0_io_dataRead : _T_386; // @[GraphicEngineVGA.scala 290:44]
  assign backBufferShadowMemories_1_clock = clock;
  assign backBufferShadowMemories_1_io_address = restoreEnabled ? _T_397 : _T_400; // @[GraphicEngineVGA.scala 287:42]
  assign backBufferShadowMemories_1_io_writeEnable = restoreEnabled ? _T_402 : _T_404; // @[GraphicEngineVGA.scala 289:46]
  assign backBufferShadowMemories_1_io_dataWrite = restoreEnabled ? backBufferRestoreMemories_1_io_dataRead : _T_406; // @[GraphicEngineVGA.scala 290:44]
  assign backBufferRestoreMemories_0_clock = clock;
  assign backBufferRestoreMemories_0_io_address = backMemoryRestoreCounter[10:0]; // @[GraphicEngineVGA.scala 282:43]
  assign backBufferRestoreMemories_1_clock = clock;
  assign backBufferRestoreMemories_1_io_address = backMemoryRestoreCounter[10:0]; // @[GraphicEngineVGA.scala 282:43]
  assign spriteMemories_0_clock = clock;
  assign spriteMemories_0_io_address = _T_537[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_1_clock = clock;
  assign spriteMemories_1_io_address = _T_656[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_2_clock = clock;
  assign spriteMemories_2_io_address = _T_775[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_3_clock = clock;
  assign spriteMemories_3_io_address = _T_894[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_4_clock = clock;
  assign spriteMemories_4_io_address = _T_1013[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_5_clock = clock;
  assign spriteMemories_5_io_address = _T_1132[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_6_clock = clock;
  assign spriteMemories_6_io_address = _T_1251[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_7_clock = clock;
  assign spriteMemories_7_io_address = _T_1370[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_8_clock = clock;
  assign spriteMemories_8_io_address = _T_1489[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_9_clock = clock;
  assign spriteMemories_9_io_address = _T_1608[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_10_clock = clock;
  assign spriteMemories_10_io_address = _T_1727[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_11_clock = clock;
  assign spriteMemories_11_io_address = _T_1846[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_12_clock = clock;
  assign spriteMemories_12_io_address = _T_1965[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_13_clock = clock;
  assign spriteMemories_13_io_address = _T_2084[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_14_clock = clock;
  assign spriteMemories_14_io_address = _T_2203[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_15_clock = clock;
  assign spriteMemories_15_io_address = _T_2322[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_16_clock = clock;
  assign spriteMemories_16_io_address = _T_2441[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_17_clock = clock;
  assign spriteMemories_17_io_address = _T_2560[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_18_clock = clock;
  assign spriteMemories_18_io_address = _T_2679[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_19_clock = clock;
  assign spriteMemories_19_io_address = _T_2798[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_20_clock = clock;
  assign spriteMemories_20_io_address = _T_2917[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_21_clock = clock;
  assign spriteMemories_21_io_address = _T_3036[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_22_clock = clock;
  assign spriteMemories_22_io_address = _T_3155[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_23_clock = clock;
  assign spriteMemories_23_io_address = _T_3274[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_24_clock = clock;
  assign spriteMemories_24_io_address = _T_3393[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_25_clock = clock;
  assign spriteMemories_25_io_address = _T_3512[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_26_clock = clock;
  assign spriteMemories_26_io_address = _T_3631[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_27_clock = clock;
  assign spriteMemories_27_io_address = _T_3750[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_28_clock = clock;
  assign spriteMemories_28_io_address = _T_3869[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_29_clock = clock;
  assign spriteMemories_29_io_address = _T_3988[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_30_clock = clock;
  assign spriteMemories_30_io_address = _T_4107[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_31_clock = clock;
  assign spriteMemories_31_io_address = _T_4226[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_32_clock = clock;
  assign spriteMemories_32_io_address = _T_4345[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_33_clock = clock;
  assign spriteMemories_33_io_address = _T_4464[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_34_clock = clock;
  assign spriteMemories_34_io_address = _T_4583[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_35_clock = clock;
  assign spriteMemories_35_io_address = _T_4702[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_36_clock = clock;
  assign spriteMemories_36_io_address = _T_4821[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_37_clock = clock;
  assign spriteMemories_37_io_address = _T_4940[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_38_clock = clock;
  assign spriteMemories_38_io_address = _T_5059[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_39_clock = clock;
  assign spriteMemories_39_io_address = _T_5178[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_40_clock = clock;
  assign spriteMemories_40_io_address = _T_5297[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_41_clock = clock;
  assign spriteMemories_41_io_address = _T_5416[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_42_clock = clock;
  assign spriteMemories_42_io_address = _T_5535[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_43_clock = clock;
  assign spriteMemories_43_io_address = _T_5654[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_44_clock = clock;
  assign spriteMemories_44_io_address = _T_5773[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_45_clock = clock;
  assign spriteMemories_45_io_address = _T_5892[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_46_clock = clock;
  assign spriteMemories_46_io_address = _T_6011[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_47_clock = clock;
  assign spriteMemories_47_io_address = _T_6130[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_48_clock = clock;
  assign spriteMemories_48_io_address = _T_6249[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_49_clock = clock;
  assign spriteMemories_49_io_address = _T_6368[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_50_clock = clock;
  assign spriteMemories_50_io_address = _T_6487[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_51_clock = clock;
  assign spriteMemories_51_io_address = _T_6606[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_52_clock = clock;
  assign spriteMemories_52_io_address = _T_6725[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_53_clock = clock;
  assign spriteMemories_53_io_address = _T_6844[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_54_clock = clock;
  assign spriteMemories_54_io_address = _T_6963[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_55_clock = clock;
  assign spriteMemories_55_io_address = _T_7082[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_56_clock = clock;
  assign spriteMemories_56_io_address = _T_7201[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_57_clock = clock;
  assign spriteMemories_57_io_address = _T_7320[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_58_clock = clock;
  assign spriteMemories_58_io_address = _T_7439[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_59_clock = clock;
  assign spriteMemories_59_io_address = _T_7558[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_60_clock = clock;
  assign spriteMemories_60_io_address = _T_7677[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_61_clock = clock;
  assign spriteMemories_61_io_address = _T_7796[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_62_clock = clock;
  assign spriteMemories_62_io_address = _T_7915[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_63_clock = clock;
  assign spriteMemories_63_io_address = _T_8034[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_64_clock = clock;
  assign spriteMemories_64_io_address = _T_8153[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_65_clock = clock;
  assign spriteMemories_65_io_address = _T_8272[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_66_clock = clock;
  assign spriteMemories_66_io_address = _T_8391[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_67_clock = clock;
  assign spriteMemories_67_io_address = _T_8510[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_68_clock = clock;
  assign spriteMemories_68_io_address = _T_8629[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_69_clock = clock;
  assign spriteMemories_69_io_address = _T_8748[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_70_clock = clock;
  assign spriteMemories_70_io_address = _T_8867[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_71_clock = clock;
  assign spriteMemories_71_io_address = _T_8986[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_72_clock = clock;
  assign spriteMemories_72_io_address = _T_9105[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_73_clock = clock;
  assign spriteMemories_73_io_address = _T_9224[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_74_clock = clock;
  assign spriteMemories_74_io_address = _T_9343[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_75_clock = clock;
  assign spriteMemories_75_io_address = _T_9462[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_76_clock = clock;
  assign spriteMemories_76_io_address = _T_9581[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_77_clock = clock;
  assign spriteMemories_77_io_address = _T_9700[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_78_clock = clock;
  assign spriteMemories_78_io_address = _T_9819[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_79_clock = clock;
  assign spriteMemories_79_io_address = _T_9938[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_80_clock = clock;
  assign spriteMemories_80_io_address = _T_10057[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_81_clock = clock;
  assign spriteMemories_81_io_address = _T_10176[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_82_clock = clock;
  assign spriteMemories_82_io_address = _T_10295[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_83_clock = clock;
  assign spriteMemories_83_io_address = _T_10414[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_84_clock = clock;
  assign spriteMemories_84_io_address = _T_10533[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_85_clock = clock;
  assign spriteMemories_85_io_address = _T_10652[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_86_clock = clock;
  assign spriteMemories_86_io_address = _T_10771[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_87_clock = clock;
  assign spriteMemories_87_io_address = _T_10890[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_88_clock = clock;
  assign spriteMemories_88_io_address = _T_11009[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_89_clock = clock;
  assign spriteMemories_89_io_address = _T_11128[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_90_clock = clock;
  assign spriteMemories_90_io_address = _T_11247[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_91_clock = clock;
  assign spriteMemories_91_io_address = _T_11366[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_92_clock = clock;
  assign spriteMemories_92_io_address = _T_11485[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_93_clock = clock;
  assign spriteMemories_93_io_address = _T_11604[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_94_clock = clock;
  assign spriteMemories_94_io_address = _T_11723[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_95_clock = clock;
  assign spriteMemories_95_io_address = _T_11842[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_96_clock = clock;
  assign spriteMemories_96_io_address = _T_11961[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_97_clock = clock;
  assign spriteMemories_97_io_address = _T_12080[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_98_clock = clock;
  assign spriteMemories_98_io_address = _T_12199[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_99_clock = clock;
  assign spriteMemories_99_io_address = _T_12318[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_100_clock = clock;
  assign spriteMemories_100_io_address = _T_12437[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_101_clock = clock;
  assign spriteMemories_101_io_address = _T_12556[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_102_clock = clock;
  assign spriteMemories_102_io_address = _T_12675[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_103_clock = clock;
  assign spriteMemories_103_io_address = _T_12794[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_104_clock = clock;
  assign spriteMemories_104_io_address = _T_12913[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_105_clock = clock;
  assign spriteMemories_105_io_address = _T_13032[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_106_clock = clock;
  assign spriteMemories_106_io_address = _T_13151[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_107_clock = clock;
  assign spriteMemories_107_io_address = _T_13270[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_108_clock = clock;
  assign spriteMemories_108_io_address = _T_13389[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_109_clock = clock;
  assign spriteMemories_109_io_address = _T_13508[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_110_clock = clock;
  assign spriteMemories_110_io_address = _T_13627[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_111_clock = clock;
  assign spriteMemories_111_io_address = _T_13746[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_112_clock = clock;
  assign spriteMemories_112_io_address = _T_13865[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_113_clock = clock;
  assign spriteMemories_113_io_address = _T_13984[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_114_clock = clock;
  assign spriteMemories_114_io_address = _T_14103[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_115_clock = clock;
  assign spriteMemories_115_io_address = _T_14222[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_116_clock = clock;
  assign spriteMemories_116_io_address = _T_14341[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_117_clock = clock;
  assign spriteMemories_117_io_address = _T_14460[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_118_clock = clock;
  assign spriteMemories_118_io_address = _T_14579[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_119_clock = clock;
  assign spriteMemories_119_io_address = _T_14698[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_120_clock = clock;
  assign spriteMemories_120_io_address = _T_14817[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_121_clock = clock;
  assign spriteMemories_121_io_address = _T_14936[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_122_clock = clock;
  assign spriteMemories_122_io_address = _T_15055[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_123_clock = clock;
  assign spriteMemories_123_io_address = _T_15174[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_124_clock = clock;
  assign spriteMemories_124_io_address = _T_15293[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_125_clock = clock;
  assign spriteMemories_125_io_address = _T_15412[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_126_clock = clock;
  assign spriteMemories_126_io_address = _T_15531[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign spriteMemories_127_clock = clock;
  assign spriteMemories_127_io_address = _T_15650[9:0]; // @[GraphicEngineVGA.scala 406:38]
  assign rotation45deg_0_clock = clock;
  assign rotation45deg_0_io_address = _T_537[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_1_clock = clock;
  assign rotation45deg_1_io_address = _T_656[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_2_clock = clock;
  assign rotation45deg_2_io_address = _T_775[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_3_clock = clock;
  assign rotation45deg_3_io_address = _T_894[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_4_clock = clock;
  assign rotation45deg_4_io_address = _T_1013[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_5_clock = clock;
  assign rotation45deg_5_io_address = _T_1132[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_6_clock = clock;
  assign rotation45deg_6_io_address = _T_1251[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_7_clock = clock;
  assign rotation45deg_7_io_address = _T_1370[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_8_clock = clock;
  assign rotation45deg_8_io_address = _T_1489[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_9_clock = clock;
  assign rotation45deg_9_io_address = _T_1608[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_10_clock = clock;
  assign rotation45deg_10_io_address = _T_1727[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_11_clock = clock;
  assign rotation45deg_11_io_address = _T_1846[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_12_clock = clock;
  assign rotation45deg_12_io_address = _T_1965[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_13_clock = clock;
  assign rotation45deg_13_io_address = _T_2084[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_14_clock = clock;
  assign rotation45deg_14_io_address = _T_2203[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_15_clock = clock;
  assign rotation45deg_15_io_address = _T_2322[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_16_clock = clock;
  assign rotation45deg_16_io_address = _T_2441[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_17_clock = clock;
  assign rotation45deg_17_io_address = _T_2560[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_18_clock = clock;
  assign rotation45deg_18_io_address = _T_2679[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_19_clock = clock;
  assign rotation45deg_19_io_address = _T_2798[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_20_clock = clock;
  assign rotation45deg_20_io_address = _T_2917[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_21_clock = clock;
  assign rotation45deg_21_io_address = _T_3036[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_22_clock = clock;
  assign rotation45deg_22_io_address = _T_3155[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_23_clock = clock;
  assign rotation45deg_23_io_address = _T_3274[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_24_clock = clock;
  assign rotation45deg_24_io_address = _T_3393[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_25_clock = clock;
  assign rotation45deg_25_io_address = _T_3512[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_26_clock = clock;
  assign rotation45deg_26_io_address = _T_3631[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_27_clock = clock;
  assign rotation45deg_27_io_address = _T_3750[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_28_clock = clock;
  assign rotation45deg_28_io_address = _T_3869[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_29_clock = clock;
  assign rotation45deg_29_io_address = _T_3988[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_30_clock = clock;
  assign rotation45deg_30_io_address = _T_4107[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_31_clock = clock;
  assign rotation45deg_31_io_address = _T_4226[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_32_clock = clock;
  assign rotation45deg_32_io_address = _T_4345[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_33_clock = clock;
  assign rotation45deg_33_io_address = _T_4464[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_34_clock = clock;
  assign rotation45deg_34_io_address = _T_4583[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_35_clock = clock;
  assign rotation45deg_35_io_address = _T_4702[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_36_clock = clock;
  assign rotation45deg_36_io_address = _T_4821[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_37_clock = clock;
  assign rotation45deg_37_io_address = _T_4940[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_38_clock = clock;
  assign rotation45deg_38_io_address = _T_5059[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_39_clock = clock;
  assign rotation45deg_39_io_address = _T_5178[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_40_clock = clock;
  assign rotation45deg_40_io_address = _T_5297[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_41_clock = clock;
  assign rotation45deg_41_io_address = _T_5416[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_42_clock = clock;
  assign rotation45deg_42_io_address = _T_5535[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_43_clock = clock;
  assign rotation45deg_43_io_address = _T_5654[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_44_clock = clock;
  assign rotation45deg_44_io_address = _T_5773[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_45_clock = clock;
  assign rotation45deg_45_io_address = _T_5892[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_46_clock = clock;
  assign rotation45deg_46_io_address = _T_6011[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_47_clock = clock;
  assign rotation45deg_47_io_address = _T_6130[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_48_clock = clock;
  assign rotation45deg_48_io_address = _T_6249[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_49_clock = clock;
  assign rotation45deg_49_io_address = _T_6368[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_50_clock = clock;
  assign rotation45deg_50_io_address = _T_6487[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_51_clock = clock;
  assign rotation45deg_51_io_address = _T_6606[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_52_clock = clock;
  assign rotation45deg_52_io_address = _T_6725[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_53_clock = clock;
  assign rotation45deg_53_io_address = _T_6844[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_54_clock = clock;
  assign rotation45deg_54_io_address = _T_6963[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_55_clock = clock;
  assign rotation45deg_55_io_address = _T_7082[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_56_clock = clock;
  assign rotation45deg_56_io_address = _T_7201[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_57_clock = clock;
  assign rotation45deg_57_io_address = _T_7320[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_58_clock = clock;
  assign rotation45deg_58_io_address = _T_7439[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_59_clock = clock;
  assign rotation45deg_59_io_address = _T_7558[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_60_clock = clock;
  assign rotation45deg_60_io_address = _T_7677[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_61_clock = clock;
  assign rotation45deg_61_io_address = _T_7796[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_62_clock = clock;
  assign rotation45deg_62_io_address = _T_7915[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_63_clock = clock;
  assign rotation45deg_63_io_address = _T_8034[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_64_clock = clock;
  assign rotation45deg_64_io_address = _T_8153[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_65_clock = clock;
  assign rotation45deg_65_io_address = _T_8272[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_66_clock = clock;
  assign rotation45deg_66_io_address = _T_8391[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_67_clock = clock;
  assign rotation45deg_67_io_address = _T_8510[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_68_clock = clock;
  assign rotation45deg_68_io_address = _T_8629[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_69_clock = clock;
  assign rotation45deg_69_io_address = _T_8748[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_70_clock = clock;
  assign rotation45deg_70_io_address = _T_8867[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_71_clock = clock;
  assign rotation45deg_71_io_address = _T_8986[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_72_clock = clock;
  assign rotation45deg_72_io_address = _T_9105[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_73_clock = clock;
  assign rotation45deg_73_io_address = _T_9224[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_74_clock = clock;
  assign rotation45deg_74_io_address = _T_9343[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_75_clock = clock;
  assign rotation45deg_75_io_address = _T_9462[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_76_clock = clock;
  assign rotation45deg_76_io_address = _T_9581[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_77_clock = clock;
  assign rotation45deg_77_io_address = _T_9700[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_78_clock = clock;
  assign rotation45deg_78_io_address = _T_9819[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_79_clock = clock;
  assign rotation45deg_79_io_address = _T_9938[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_80_clock = clock;
  assign rotation45deg_80_io_address = _T_10057[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_81_clock = clock;
  assign rotation45deg_81_io_address = _T_10176[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_82_clock = clock;
  assign rotation45deg_82_io_address = _T_10295[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_83_clock = clock;
  assign rotation45deg_83_io_address = _T_10414[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_84_clock = clock;
  assign rotation45deg_84_io_address = _T_10533[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_85_clock = clock;
  assign rotation45deg_85_io_address = _T_10652[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_86_clock = clock;
  assign rotation45deg_86_io_address = _T_10771[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_87_clock = clock;
  assign rotation45deg_87_io_address = _T_10890[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_88_clock = clock;
  assign rotation45deg_88_io_address = _T_11009[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_89_clock = clock;
  assign rotation45deg_89_io_address = _T_11128[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_90_clock = clock;
  assign rotation45deg_90_io_address = _T_11247[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_91_clock = clock;
  assign rotation45deg_91_io_address = _T_11366[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_92_clock = clock;
  assign rotation45deg_92_io_address = _T_11485[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_93_clock = clock;
  assign rotation45deg_93_io_address = _T_11604[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_94_clock = clock;
  assign rotation45deg_94_io_address = _T_11723[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_95_clock = clock;
  assign rotation45deg_95_io_address = _T_11842[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_96_clock = clock;
  assign rotation45deg_96_io_address = _T_11961[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_97_clock = clock;
  assign rotation45deg_97_io_address = _T_12080[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_98_clock = clock;
  assign rotation45deg_98_io_address = _T_12199[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_99_clock = clock;
  assign rotation45deg_99_io_address = _T_12318[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_100_clock = clock;
  assign rotation45deg_100_io_address = _T_12437[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_101_clock = clock;
  assign rotation45deg_101_io_address = _T_12556[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_102_clock = clock;
  assign rotation45deg_102_io_address = _T_12675[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_103_clock = clock;
  assign rotation45deg_103_io_address = _T_12794[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_104_clock = clock;
  assign rotation45deg_104_io_address = _T_12913[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_105_clock = clock;
  assign rotation45deg_105_io_address = _T_13032[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_106_clock = clock;
  assign rotation45deg_106_io_address = _T_13151[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_107_clock = clock;
  assign rotation45deg_107_io_address = _T_13270[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_108_clock = clock;
  assign rotation45deg_108_io_address = _T_13389[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_109_clock = clock;
  assign rotation45deg_109_io_address = _T_13508[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_110_clock = clock;
  assign rotation45deg_110_io_address = _T_13627[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_111_clock = clock;
  assign rotation45deg_111_io_address = _T_13746[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_112_clock = clock;
  assign rotation45deg_112_io_address = _T_13865[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_113_clock = clock;
  assign rotation45deg_113_io_address = _T_13984[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_114_clock = clock;
  assign rotation45deg_114_io_address = _T_14103[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_115_clock = clock;
  assign rotation45deg_115_io_address = _T_14222[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_116_clock = clock;
  assign rotation45deg_116_io_address = _T_14341[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_117_clock = clock;
  assign rotation45deg_117_io_address = _T_14460[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_118_clock = clock;
  assign rotation45deg_118_io_address = _T_14579[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_119_clock = clock;
  assign rotation45deg_119_io_address = _T_14698[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_120_clock = clock;
  assign rotation45deg_120_io_address = _T_14817[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_121_clock = clock;
  assign rotation45deg_121_io_address = _T_14936[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_122_clock = clock;
  assign rotation45deg_122_io_address = _T_15055[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_123_clock = clock;
  assign rotation45deg_123_io_address = _T_15174[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_124_clock = clock;
  assign rotation45deg_124_io_address = _T_15293[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_125_clock = clock;
  assign rotation45deg_125_io_address = _T_15412[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_126_clock = clock;
  assign rotation45deg_126_io_address = _T_15531[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign rotation45deg_127_clock = clock;
  assign rotation45deg_127_io_address = _T_15650[11:0]; // @[GraphicEngineVGA.scala 402:33]
  assign spriteBlender_clock = clock;
  assign spriteBlender_io_pixelColorBack = pixelColorBack; // @[GraphicEngineVGA.scala 337:35]
  assign spriteBlender_io_spriteVisibleReg_0 = spriteVisibleReg_0; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_1 = spriteVisibleReg_1; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_2 = spriteVisibleReg_2; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_3 = spriteVisibleReg_3; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_4 = spriteVisibleReg_4; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_5 = spriteVisibleReg_5; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_6 = spriteVisibleReg_6; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_7 = spriteVisibleReg_7; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_8 = spriteVisibleReg_8; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_9 = spriteVisibleReg_9; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_10 = spriteVisibleReg_10; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_11 = spriteVisibleReg_11; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_12 = spriteVisibleReg_12; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_13 = spriteVisibleReg_13; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_14 = spriteVisibleReg_14; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_15 = spriteVisibleReg_15; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_16 = spriteVisibleReg_16; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_17 = spriteVisibleReg_17; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_18 = spriteVisibleReg_18; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_19 = spriteVisibleReg_19; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_20 = spriteVisibleReg_20; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_21 = spriteVisibleReg_21; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_22 = spriteVisibleReg_22; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_23 = spriteVisibleReg_23; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_24 = spriteVisibleReg_24; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_25 = spriteVisibleReg_25; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_26 = spriteVisibleReg_26; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_27 = spriteVisibleReg_27; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_28 = spriteVisibleReg_28; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_29 = spriteVisibleReg_29; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_30 = spriteVisibleReg_30; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_31 = spriteVisibleReg_31; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_32 = spriteVisibleReg_32; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_33 = spriteVisibleReg_33; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_41 = spriteVisibleReg_41; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_42 = spriteVisibleReg_42; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_43 = spriteVisibleReg_43; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_44 = spriteVisibleReg_44; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_45 = spriteVisibleReg_45; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_46 = spriteVisibleReg_46; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_47 = spriteVisibleReg_47; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_48 = spriteVisibleReg_48; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_49 = spriteVisibleReg_49; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_50 = spriteVisibleReg_50; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_51 = spriteVisibleReg_51; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_55 = spriteVisibleReg_55; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_56 = spriteVisibleReg_56; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_57 = spriteVisibleReg_57; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_61 = spriteVisibleReg_61; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_62 = spriteVisibleReg_62; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_63 = spriteVisibleReg_63; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_64 = spriteVisibleReg_64; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_65 = spriteVisibleReg_65; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_66 = spriteVisibleReg_66; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_70 = spriteVisibleReg_70; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_71 = spriteVisibleReg_71; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_spriteVisibleReg_72 = spriteVisibleReg_72; // @[GraphicEngineVGA.scala 338:37]
  assign spriteBlender_io_inSprite_0 = _T_509 & _T_512; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_1 = _T_628 & _T_631; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_2 = _T_747 & _T_750; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_3 = _T_866 & _T_869; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_4 = _T_985 & _T_988; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_5 = _T_1104 & _T_1107; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_6 = _T_1223 & _T_1226; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_7 = _T_1342 & _T_1345; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_8 = _T_1461 & _T_1464; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_9 = _T_1580 & _T_1583; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_10 = _T_1699 & _T_1702; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_11 = _T_1818 & _T_1821; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_12 = _T_1937 & _T_1940; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_13 = _T_2056 & _T_2059; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_14 = _T_2175 & _T_2178; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_15 = _T_2294 & _T_2297; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_16 = _T_2413 & _T_2416; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_17 = _T_2532 & _T_2535; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_18 = _T_2651 & _T_2654; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_19 = _T_2770 & _T_2773; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_20 = _T_2889 & _T_2892; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_21 = _T_3008 & _T_3011; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_22 = _T_3127 & _T_3130; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_23 = _T_3246 & _T_3249; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_24 = _T_3365 & _T_3368; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_25 = _T_3484 & _T_3487; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_26 = _T_3603 & _T_3606; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_27 = _T_3722 & _T_3725; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_28 = _T_3841 & _T_3844; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_29 = _T_3960 & _T_3963; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_30 = _T_4079 & _T_4082; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_31 = _T_4198 & _T_4201; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_32 = _T_4317 & _T_4320; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_33 = _T_4436 & _T_4439; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_34 = _T_4555 & _T_4558; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_35 = _T_4674 & _T_4677; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_36 = _T_4793 & _T_4796; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_37 = _T_4912 & _T_4915; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_38 = _T_5031 & _T_5034; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_39 = _T_5150 & _T_5153; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_40 = _T_5269 & _T_5272; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_41 = _T_5388 & _T_5391; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_42 = _T_5507 & _T_5510; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_43 = _T_5626 & _T_5629; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_44 = _T_5745 & _T_5748; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_45 = _T_5864 & _T_5867; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_46 = _T_5983 & _T_5986; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_47 = _T_6102 & _T_6105; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_48 = _T_6221 & _T_6224; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_49 = _T_6340 & _T_6343; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_50 = _T_6459 & _T_6462; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_51 = _T_6578 & _T_6581; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_52 = _T_6697 & _T_6700; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_53 = _T_6816 & _T_6819; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_54 = _T_6935 & _T_6938; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_55 = _T_7054 & _T_7057; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_56 = _T_7173 & _T_7176; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_57 = _T_7292 & _T_7295; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_58 = _T_7411 & _T_7414; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_59 = _T_7530 & _T_7533; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_60 = _T_7649 & _T_7652; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_61 = _T_7768 & _T_7771; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_62 = _T_7887 & _T_7890; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_63 = _T_8006 & _T_8009; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_64 = _T_8125 & _T_8128; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_65 = _T_8244 & _T_8247; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_66 = _T_8363 & _T_8366; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_67 = _T_8482 & _T_8485; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_68 = _T_8601 & _T_8604; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_69 = _T_8720 & _T_8723; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_70 = _T_8839 & _T_8842; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_71 = _T_8958 & _T_8961; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_72 = _T_9077 & _T_9080; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_73 = _T_9196 & _T_9199; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_74 = _T_9315 & _T_9318; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_75 = _T_9434 & _T_9437; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_76 = _T_9553 & _T_9556; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_77 = _T_9672 & _T_9675; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_78 = _T_9791 & _T_9794; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_79 = _T_9910 & _T_9913; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_80 = _T_10029 & _T_10032; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_81 = _T_10148 & _T_10151; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_82 = _T_10267 & _T_10270; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_83 = _T_10386 & _T_10389; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_84 = _T_10505 & _T_10508; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_85 = _T_10624 & _T_10627; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_86 = _T_10743 & _T_10746; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_87 = _T_10862 & _T_10865; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_88 = _T_10981 & _T_10984; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_89 = _T_11100 & _T_11103; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_90 = _T_11219 & _T_11222; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_91 = _T_11338 & _T_11341; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_92 = _T_11457 & _T_11460; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_93 = _T_11576 & _T_11579; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_94 = _T_11695 & _T_11698; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_95 = _T_11814 & _T_11817; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_96 = _T_11933 & _T_11936; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_97 = _T_12052 & _T_12055; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_98 = _T_12171 & _T_12174; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_99 = _T_12290 & _T_12293; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_100 = _T_12409 & _T_12412; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_101 = _T_12528 & _T_12531; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_102 = _T_12647 & _T_12650; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_103 = _T_12766 & _T_12769; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_104 = _T_12885 & _T_12888; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_105 = _T_13004 & _T_13007; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_106 = _T_13123 & _T_13126; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_107 = _T_13242 & _T_13245; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_108 = _T_13361 & _T_13364; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_109 = _T_13480 & _T_13483; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_110 = _T_13599 & _T_13602; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_111 = _T_13718 & _T_13721; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_112 = _T_13837 & _T_13840; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_113 = _T_13956 & _T_13959; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_114 = _T_14075 & _T_14078; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_115 = _T_14194 & _T_14197; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_116 = _T_14313 & _T_14316; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_117 = _T_14432 & _T_14435; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_118 = _T_14551 & _T_14554; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_119 = _T_14670 & _T_14673; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_120 = _T_14789 & _T_14792; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_121 = _T_14908 & _T_14911; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_122 = _T_15027 & _T_15030; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_123 = _T_15146 & _T_15149; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_124 = _T_15265 & _T_15268; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_125 = _T_15384 & _T_15387; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_126 = _T_15503 & _T_15506; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_inSprite_127 = _T_15622 & _T_15625; // @[GraphicEngineVGA.scala 339:28]
  assign spriteBlender_io_datareader_0 = spriteMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_1 = spriteMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_2 = spriteMemories_2_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_3 = spriteMemories_3_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_4 = spriteMemories_4_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_5 = spriteMemories_5_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_6 = spriteMemories_6_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_7 = spriteMemories_7_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_8 = spriteMemories_8_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_9 = spriteMemories_9_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_10 = spriteMemories_10_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_11 = spriteMemories_11_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_12 = spriteMemories_12_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_13 = spriteMemories_13_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_14 = spriteMemories_14_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_15 = spriteMemories_15_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_16 = spriteMemories_16_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_17 = spriteMemories_17_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_18 = spriteMemories_18_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_19 = spriteMemories_19_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_20 = spriteMemories_20_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_21 = spriteMemories_21_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_22 = spriteMemories_22_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_23 = spriteMemories_23_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_24 = spriteMemories_24_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_25 = spriteMemories_25_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_26 = spriteMemories_26_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_27 = spriteMemories_27_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_28 = spriteMemories_28_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_29 = spriteMemories_29_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_30 = spriteMemories_30_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_31 = spriteMemories_31_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_32 = spriteMemories_32_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_33 = spriteMemories_33_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_34 = spriteMemories_34_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_35 = spriteMemories_35_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_36 = spriteMemories_36_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_37 = spriteMemories_37_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_38 = spriteMemories_38_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_39 = spriteMemories_39_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_40 = spriteMemories_40_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_41 = spriteMemories_41_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_42 = spriteMemories_42_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_43 = spriteMemories_43_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_44 = spriteMemories_44_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_45 = spriteMemories_45_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_46 = spriteMemories_46_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_47 = spriteMemories_47_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_48 = spriteMemories_48_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_49 = spriteMemories_49_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_50 = spriteMemories_50_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_51 = spriteMemories_51_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_52 = spriteMemories_52_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_53 = spriteMemories_53_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_54 = spriteMemories_54_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_55 = spriteMemories_55_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_56 = spriteMemories_56_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_57 = spriteMemories_57_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_58 = spriteMemories_58_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_59 = spriteMemories_59_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_60 = spriteMemories_60_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_61 = spriteMemories_61_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_62 = spriteMemories_62_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_63 = spriteMemories_63_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_64 = spriteMemories_64_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_65 = spriteMemories_65_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_66 = spriteMemories_66_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_67 = spriteMemories_67_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_68 = spriteMemories_68_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_69 = spriteMemories_69_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_70 = spriteMemories_70_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_71 = spriteMemories_71_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_72 = spriteMemories_72_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_73 = spriteMemories_73_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_74 = spriteMemories_74_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_75 = spriteMemories_75_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_76 = spriteMemories_76_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_77 = spriteMemories_77_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_78 = spriteMemories_78_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_79 = spriteMemories_79_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_80 = spriteMemories_80_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_81 = spriteMemories_81_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_82 = spriteMemories_82_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_83 = spriteMemories_83_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_84 = spriteMemories_84_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_85 = spriteMemories_85_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_86 = spriteMemories_86_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_87 = spriteMemories_87_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_88 = spriteMemories_88_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_89 = spriteMemories_89_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_90 = spriteMemories_90_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_91 = spriteMemories_91_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_92 = spriteMemories_92_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_93 = spriteMemories_93_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_94 = spriteMemories_94_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_95 = spriteMemories_95_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_96 = spriteMemories_96_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_97 = spriteMemories_97_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_98 = spriteMemories_98_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_99 = spriteMemories_99_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_100 = spriteMemories_100_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_101 = spriteMemories_101_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_102 = spriteMemories_102_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_103 = spriteMemories_103_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_104 = spriteMemories_104_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_105 = spriteMemories_105_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_106 = spriteMemories_106_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_107 = spriteMemories_107_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_108 = spriteMemories_108_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_109 = spriteMemories_109_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_110 = spriteMemories_110_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_111 = spriteMemories_111_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_112 = spriteMemories_112_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_113 = spriteMemories_113_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_114 = spriteMemories_114_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_115 = spriteMemories_115_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_116 = spriteMemories_116_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_117 = spriteMemories_117_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_118 = spriteMemories_118_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_119 = spriteMemories_119_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_120 = spriteMemories_120_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_121 = spriteMemories_121_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_122 = spriteMemories_122_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_123 = spriteMemories_123_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_124 = spriteMemories_124_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_125 = spriteMemories_125_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_126 = spriteMemories_126_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
  assign spriteBlender_io_datareader_127 = spriteMemories_127_io_dataRead; // @[GraphicEngineVGA.scala 407:36]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ScaleCounterReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  CounterXReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  CounterYReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  backMemoryRestoreCounter = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  _T_14_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_14_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_14_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_14_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_16_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_16_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_16_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_16_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  frameClockCount = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXPositionReg_0 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXPositionReg_1 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXPositionReg_2 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXPositionReg_3 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXPositionReg_4 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXPositionReg_5 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXPositionReg_6 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXPositionReg_7 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXPositionReg_8 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXPositionReg_9 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXPositionReg_10 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXPositionReg_11 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXPositionReg_12 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXPositionReg_13 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXPositionReg_14 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXPositionReg_15 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXPositionReg_16 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXPositionReg_17 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXPositionReg_18 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXPositionReg_19 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXPositionReg_20 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXPositionReg_21 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXPositionReg_22 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXPositionReg_23 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXPositionReg_24 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXPositionReg_25 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXPositionReg_26 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXPositionReg_27 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXPositionReg_28 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXPositionReg_29 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXPositionReg_30 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXPositionReg_31 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXPositionReg_32 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXPositionReg_33 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXPositionReg_34 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXPositionReg_35 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXPositionReg_36 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXPositionReg_37 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXPositionReg_38 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXPositionReg_39 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXPositionReg_40 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXPositionReg_41 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXPositionReg_42 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXPositionReg_43 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXPositionReg_44 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteXPositionReg_45 = _RAND_58[10:0];
  _RAND_59 = {1{`RANDOM}};
  spriteXPositionReg_46 = _RAND_59[10:0];
  _RAND_60 = {1{`RANDOM}};
  spriteXPositionReg_47 = _RAND_60[10:0];
  _RAND_61 = {1{`RANDOM}};
  spriteXPositionReg_48 = _RAND_61[10:0];
  _RAND_62 = {1{`RANDOM}};
  spriteXPositionReg_49 = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  spriteXPositionReg_50 = _RAND_63[10:0];
  _RAND_64 = {1{`RANDOM}};
  spriteXPositionReg_51 = _RAND_64[10:0];
  _RAND_65 = {1{`RANDOM}};
  spriteXPositionReg_52 = _RAND_65[10:0];
  _RAND_66 = {1{`RANDOM}};
  spriteXPositionReg_53 = _RAND_66[10:0];
  _RAND_67 = {1{`RANDOM}};
  spriteXPositionReg_54 = _RAND_67[10:0];
  _RAND_68 = {1{`RANDOM}};
  spriteXPositionReg_55 = _RAND_68[10:0];
  _RAND_69 = {1{`RANDOM}};
  spriteXPositionReg_56 = _RAND_69[10:0];
  _RAND_70 = {1{`RANDOM}};
  spriteXPositionReg_57 = _RAND_70[10:0];
  _RAND_71 = {1{`RANDOM}};
  spriteXPositionReg_58 = _RAND_71[10:0];
  _RAND_72 = {1{`RANDOM}};
  spriteXPositionReg_59 = _RAND_72[10:0];
  _RAND_73 = {1{`RANDOM}};
  spriteXPositionReg_60 = _RAND_73[10:0];
  _RAND_74 = {1{`RANDOM}};
  spriteXPositionReg_61 = _RAND_74[10:0];
  _RAND_75 = {1{`RANDOM}};
  spriteXPositionReg_62 = _RAND_75[10:0];
  _RAND_76 = {1{`RANDOM}};
  spriteXPositionReg_63 = _RAND_76[10:0];
  _RAND_77 = {1{`RANDOM}};
  spriteXPositionReg_64 = _RAND_77[10:0];
  _RAND_78 = {1{`RANDOM}};
  spriteXPositionReg_65 = _RAND_78[10:0];
  _RAND_79 = {1{`RANDOM}};
  spriteXPositionReg_66 = _RAND_79[10:0];
  _RAND_80 = {1{`RANDOM}};
  spriteXPositionReg_67 = _RAND_80[10:0];
  _RAND_81 = {1{`RANDOM}};
  spriteXPositionReg_68 = _RAND_81[10:0];
  _RAND_82 = {1{`RANDOM}};
  spriteXPositionReg_69 = _RAND_82[10:0];
  _RAND_83 = {1{`RANDOM}};
  spriteXPositionReg_70 = _RAND_83[10:0];
  _RAND_84 = {1{`RANDOM}};
  spriteXPositionReg_71 = _RAND_84[10:0];
  _RAND_85 = {1{`RANDOM}};
  spriteXPositionReg_72 = _RAND_85[10:0];
  _RAND_86 = {1{`RANDOM}};
  spriteXPositionReg_73 = _RAND_86[10:0];
  _RAND_87 = {1{`RANDOM}};
  spriteXPositionReg_74 = _RAND_87[10:0];
  _RAND_88 = {1{`RANDOM}};
  spriteXPositionReg_75 = _RAND_88[10:0];
  _RAND_89 = {1{`RANDOM}};
  spriteXPositionReg_76 = _RAND_89[10:0];
  _RAND_90 = {1{`RANDOM}};
  spriteXPositionReg_77 = _RAND_90[10:0];
  _RAND_91 = {1{`RANDOM}};
  spriteXPositionReg_78 = _RAND_91[10:0];
  _RAND_92 = {1{`RANDOM}};
  spriteXPositionReg_79 = _RAND_92[10:0];
  _RAND_93 = {1{`RANDOM}};
  spriteXPositionReg_80 = _RAND_93[10:0];
  _RAND_94 = {1{`RANDOM}};
  spriteXPositionReg_81 = _RAND_94[10:0];
  _RAND_95 = {1{`RANDOM}};
  spriteXPositionReg_82 = _RAND_95[10:0];
  _RAND_96 = {1{`RANDOM}};
  spriteXPositionReg_83 = _RAND_96[10:0];
  _RAND_97 = {1{`RANDOM}};
  spriteXPositionReg_84 = _RAND_97[10:0];
  _RAND_98 = {1{`RANDOM}};
  spriteXPositionReg_85 = _RAND_98[10:0];
  _RAND_99 = {1{`RANDOM}};
  spriteXPositionReg_86 = _RAND_99[10:0];
  _RAND_100 = {1{`RANDOM}};
  spriteXPositionReg_87 = _RAND_100[10:0];
  _RAND_101 = {1{`RANDOM}};
  spriteXPositionReg_88 = _RAND_101[10:0];
  _RAND_102 = {1{`RANDOM}};
  spriteXPositionReg_89 = _RAND_102[10:0];
  _RAND_103 = {1{`RANDOM}};
  spriteXPositionReg_90 = _RAND_103[10:0];
  _RAND_104 = {1{`RANDOM}};
  spriteXPositionReg_91 = _RAND_104[10:0];
  _RAND_105 = {1{`RANDOM}};
  spriteXPositionReg_92 = _RAND_105[10:0];
  _RAND_106 = {1{`RANDOM}};
  spriteXPositionReg_93 = _RAND_106[10:0];
  _RAND_107 = {1{`RANDOM}};
  spriteXPositionReg_94 = _RAND_107[10:0];
  _RAND_108 = {1{`RANDOM}};
  spriteXPositionReg_95 = _RAND_108[10:0];
  _RAND_109 = {1{`RANDOM}};
  spriteXPositionReg_96 = _RAND_109[10:0];
  _RAND_110 = {1{`RANDOM}};
  spriteXPositionReg_97 = _RAND_110[10:0];
  _RAND_111 = {1{`RANDOM}};
  spriteXPositionReg_98 = _RAND_111[10:0];
  _RAND_112 = {1{`RANDOM}};
  spriteXPositionReg_99 = _RAND_112[10:0];
  _RAND_113 = {1{`RANDOM}};
  spriteXPositionReg_100 = _RAND_113[10:0];
  _RAND_114 = {1{`RANDOM}};
  spriteXPositionReg_101 = _RAND_114[10:0];
  _RAND_115 = {1{`RANDOM}};
  spriteXPositionReg_102 = _RAND_115[10:0];
  _RAND_116 = {1{`RANDOM}};
  spriteXPositionReg_103 = _RAND_116[10:0];
  _RAND_117 = {1{`RANDOM}};
  spriteXPositionReg_104 = _RAND_117[10:0];
  _RAND_118 = {1{`RANDOM}};
  spriteXPositionReg_105 = _RAND_118[10:0];
  _RAND_119 = {1{`RANDOM}};
  spriteXPositionReg_106 = _RAND_119[10:0];
  _RAND_120 = {1{`RANDOM}};
  spriteXPositionReg_107 = _RAND_120[10:0];
  _RAND_121 = {1{`RANDOM}};
  spriteXPositionReg_108 = _RAND_121[10:0];
  _RAND_122 = {1{`RANDOM}};
  spriteXPositionReg_109 = _RAND_122[10:0];
  _RAND_123 = {1{`RANDOM}};
  spriteXPositionReg_110 = _RAND_123[10:0];
  _RAND_124 = {1{`RANDOM}};
  spriteXPositionReg_111 = _RAND_124[10:0];
  _RAND_125 = {1{`RANDOM}};
  spriteXPositionReg_112 = _RAND_125[10:0];
  _RAND_126 = {1{`RANDOM}};
  spriteXPositionReg_113 = _RAND_126[10:0];
  _RAND_127 = {1{`RANDOM}};
  spriteXPositionReg_114 = _RAND_127[10:0];
  _RAND_128 = {1{`RANDOM}};
  spriteXPositionReg_115 = _RAND_128[10:0];
  _RAND_129 = {1{`RANDOM}};
  spriteXPositionReg_116 = _RAND_129[10:0];
  _RAND_130 = {1{`RANDOM}};
  spriteXPositionReg_117 = _RAND_130[10:0];
  _RAND_131 = {1{`RANDOM}};
  spriteXPositionReg_118 = _RAND_131[10:0];
  _RAND_132 = {1{`RANDOM}};
  spriteXPositionReg_119 = _RAND_132[10:0];
  _RAND_133 = {1{`RANDOM}};
  spriteXPositionReg_120 = _RAND_133[10:0];
  _RAND_134 = {1{`RANDOM}};
  spriteXPositionReg_121 = _RAND_134[10:0];
  _RAND_135 = {1{`RANDOM}};
  spriteXPositionReg_122 = _RAND_135[10:0];
  _RAND_136 = {1{`RANDOM}};
  spriteXPositionReg_123 = _RAND_136[10:0];
  _RAND_137 = {1{`RANDOM}};
  spriteXPositionReg_124 = _RAND_137[10:0];
  _RAND_138 = {1{`RANDOM}};
  spriteXPositionReg_125 = _RAND_138[10:0];
  _RAND_139 = {1{`RANDOM}};
  spriteXPositionReg_126 = _RAND_139[10:0];
  _RAND_140 = {1{`RANDOM}};
  spriteXPositionReg_127 = _RAND_140[10:0];
  _RAND_141 = {1{`RANDOM}};
  spriteYPositionReg_0 = _RAND_141[9:0];
  _RAND_142 = {1{`RANDOM}};
  spriteYPositionReg_1 = _RAND_142[9:0];
  _RAND_143 = {1{`RANDOM}};
  spriteYPositionReg_2 = _RAND_143[9:0];
  _RAND_144 = {1{`RANDOM}};
  spriteYPositionReg_3 = _RAND_144[9:0];
  _RAND_145 = {1{`RANDOM}};
  spriteYPositionReg_4 = _RAND_145[9:0];
  _RAND_146 = {1{`RANDOM}};
  spriteYPositionReg_5 = _RAND_146[9:0];
  _RAND_147 = {1{`RANDOM}};
  spriteYPositionReg_6 = _RAND_147[9:0];
  _RAND_148 = {1{`RANDOM}};
  spriteYPositionReg_7 = _RAND_148[9:0];
  _RAND_149 = {1{`RANDOM}};
  spriteYPositionReg_8 = _RAND_149[9:0];
  _RAND_150 = {1{`RANDOM}};
  spriteYPositionReg_9 = _RAND_150[9:0];
  _RAND_151 = {1{`RANDOM}};
  spriteYPositionReg_10 = _RAND_151[9:0];
  _RAND_152 = {1{`RANDOM}};
  spriteYPositionReg_11 = _RAND_152[9:0];
  _RAND_153 = {1{`RANDOM}};
  spriteYPositionReg_12 = _RAND_153[9:0];
  _RAND_154 = {1{`RANDOM}};
  spriteYPositionReg_13 = _RAND_154[9:0];
  _RAND_155 = {1{`RANDOM}};
  spriteYPositionReg_14 = _RAND_155[9:0];
  _RAND_156 = {1{`RANDOM}};
  spriteYPositionReg_15 = _RAND_156[9:0];
  _RAND_157 = {1{`RANDOM}};
  spriteYPositionReg_16 = _RAND_157[9:0];
  _RAND_158 = {1{`RANDOM}};
  spriteYPositionReg_17 = _RAND_158[9:0];
  _RAND_159 = {1{`RANDOM}};
  spriteYPositionReg_18 = _RAND_159[9:0];
  _RAND_160 = {1{`RANDOM}};
  spriteYPositionReg_19 = _RAND_160[9:0];
  _RAND_161 = {1{`RANDOM}};
  spriteYPositionReg_20 = _RAND_161[9:0];
  _RAND_162 = {1{`RANDOM}};
  spriteYPositionReg_21 = _RAND_162[9:0];
  _RAND_163 = {1{`RANDOM}};
  spriteYPositionReg_22 = _RAND_163[9:0];
  _RAND_164 = {1{`RANDOM}};
  spriteYPositionReg_23 = _RAND_164[9:0];
  _RAND_165 = {1{`RANDOM}};
  spriteYPositionReg_24 = _RAND_165[9:0];
  _RAND_166 = {1{`RANDOM}};
  spriteYPositionReg_25 = _RAND_166[9:0];
  _RAND_167 = {1{`RANDOM}};
  spriteYPositionReg_26 = _RAND_167[9:0];
  _RAND_168 = {1{`RANDOM}};
  spriteYPositionReg_27 = _RAND_168[9:0];
  _RAND_169 = {1{`RANDOM}};
  spriteYPositionReg_28 = _RAND_169[9:0];
  _RAND_170 = {1{`RANDOM}};
  spriteYPositionReg_29 = _RAND_170[9:0];
  _RAND_171 = {1{`RANDOM}};
  spriteYPositionReg_30 = _RAND_171[9:0];
  _RAND_172 = {1{`RANDOM}};
  spriteYPositionReg_31 = _RAND_172[9:0];
  _RAND_173 = {1{`RANDOM}};
  spriteYPositionReg_32 = _RAND_173[9:0];
  _RAND_174 = {1{`RANDOM}};
  spriteYPositionReg_33 = _RAND_174[9:0];
  _RAND_175 = {1{`RANDOM}};
  spriteYPositionReg_34 = _RAND_175[9:0];
  _RAND_176 = {1{`RANDOM}};
  spriteYPositionReg_35 = _RAND_176[9:0];
  _RAND_177 = {1{`RANDOM}};
  spriteYPositionReg_36 = _RAND_177[9:0];
  _RAND_178 = {1{`RANDOM}};
  spriteYPositionReg_37 = _RAND_178[9:0];
  _RAND_179 = {1{`RANDOM}};
  spriteYPositionReg_38 = _RAND_179[9:0];
  _RAND_180 = {1{`RANDOM}};
  spriteYPositionReg_39 = _RAND_180[9:0];
  _RAND_181 = {1{`RANDOM}};
  spriteYPositionReg_40 = _RAND_181[9:0];
  _RAND_182 = {1{`RANDOM}};
  spriteYPositionReg_41 = _RAND_182[9:0];
  _RAND_183 = {1{`RANDOM}};
  spriteYPositionReg_42 = _RAND_183[9:0];
  _RAND_184 = {1{`RANDOM}};
  spriteYPositionReg_43 = _RAND_184[9:0];
  _RAND_185 = {1{`RANDOM}};
  spriteYPositionReg_44 = _RAND_185[9:0];
  _RAND_186 = {1{`RANDOM}};
  spriteYPositionReg_45 = _RAND_186[9:0];
  _RAND_187 = {1{`RANDOM}};
  spriteYPositionReg_46 = _RAND_187[9:0];
  _RAND_188 = {1{`RANDOM}};
  spriteYPositionReg_47 = _RAND_188[9:0];
  _RAND_189 = {1{`RANDOM}};
  spriteYPositionReg_48 = _RAND_189[9:0];
  _RAND_190 = {1{`RANDOM}};
  spriteYPositionReg_49 = _RAND_190[9:0];
  _RAND_191 = {1{`RANDOM}};
  spriteYPositionReg_50 = _RAND_191[9:0];
  _RAND_192 = {1{`RANDOM}};
  spriteYPositionReg_51 = _RAND_192[9:0];
  _RAND_193 = {1{`RANDOM}};
  spriteYPositionReg_52 = _RAND_193[9:0];
  _RAND_194 = {1{`RANDOM}};
  spriteYPositionReg_53 = _RAND_194[9:0];
  _RAND_195 = {1{`RANDOM}};
  spriteYPositionReg_54 = _RAND_195[9:0];
  _RAND_196 = {1{`RANDOM}};
  spriteYPositionReg_55 = _RAND_196[9:0];
  _RAND_197 = {1{`RANDOM}};
  spriteYPositionReg_56 = _RAND_197[9:0];
  _RAND_198 = {1{`RANDOM}};
  spriteYPositionReg_57 = _RAND_198[9:0];
  _RAND_199 = {1{`RANDOM}};
  spriteYPositionReg_58 = _RAND_199[9:0];
  _RAND_200 = {1{`RANDOM}};
  spriteYPositionReg_59 = _RAND_200[9:0];
  _RAND_201 = {1{`RANDOM}};
  spriteYPositionReg_60 = _RAND_201[9:0];
  _RAND_202 = {1{`RANDOM}};
  spriteYPositionReg_61 = _RAND_202[9:0];
  _RAND_203 = {1{`RANDOM}};
  spriteYPositionReg_62 = _RAND_203[9:0];
  _RAND_204 = {1{`RANDOM}};
  spriteYPositionReg_63 = _RAND_204[9:0];
  _RAND_205 = {1{`RANDOM}};
  spriteYPositionReg_70 = _RAND_205[9:0];
  _RAND_206 = {1{`RANDOM}};
  spriteYPositionReg_71 = _RAND_206[9:0];
  _RAND_207 = {1{`RANDOM}};
  spriteYPositionReg_72 = _RAND_207[9:0];
  _RAND_208 = {1{`RANDOM}};
  spriteYPositionReg_73 = _RAND_208[9:0];
  _RAND_209 = {1{`RANDOM}};
  spriteYPositionReg_74 = _RAND_209[9:0];
  _RAND_210 = {1{`RANDOM}};
  spriteYPositionReg_75 = _RAND_210[9:0];
  _RAND_211 = {1{`RANDOM}};
  spriteYPositionReg_76 = _RAND_211[9:0];
  _RAND_212 = {1{`RANDOM}};
  spriteYPositionReg_77 = _RAND_212[9:0];
  _RAND_213 = {1{`RANDOM}};
  spriteYPositionReg_78 = _RAND_213[9:0];
  _RAND_214 = {1{`RANDOM}};
  spriteYPositionReg_79 = _RAND_214[9:0];
  _RAND_215 = {1{`RANDOM}};
  spriteYPositionReg_80 = _RAND_215[9:0];
  _RAND_216 = {1{`RANDOM}};
  spriteYPositionReg_81 = _RAND_216[9:0];
  _RAND_217 = {1{`RANDOM}};
  spriteYPositionReg_82 = _RAND_217[9:0];
  _RAND_218 = {1{`RANDOM}};
  spriteYPositionReg_83 = _RAND_218[9:0];
  _RAND_219 = {1{`RANDOM}};
  spriteYPositionReg_84 = _RAND_219[9:0];
  _RAND_220 = {1{`RANDOM}};
  spriteYPositionReg_85 = _RAND_220[9:0];
  _RAND_221 = {1{`RANDOM}};
  spriteYPositionReg_86 = _RAND_221[9:0];
  _RAND_222 = {1{`RANDOM}};
  spriteYPositionReg_87 = _RAND_222[9:0];
  _RAND_223 = {1{`RANDOM}};
  spriteYPositionReg_88 = _RAND_223[9:0];
  _RAND_224 = {1{`RANDOM}};
  spriteYPositionReg_89 = _RAND_224[9:0];
  _RAND_225 = {1{`RANDOM}};
  spriteYPositionReg_90 = _RAND_225[9:0];
  _RAND_226 = {1{`RANDOM}};
  spriteYPositionReg_91 = _RAND_226[9:0];
  _RAND_227 = {1{`RANDOM}};
  spriteYPositionReg_92 = _RAND_227[9:0];
  _RAND_228 = {1{`RANDOM}};
  spriteYPositionReg_93 = _RAND_228[9:0];
  _RAND_229 = {1{`RANDOM}};
  spriteYPositionReg_94 = _RAND_229[9:0];
  _RAND_230 = {1{`RANDOM}};
  spriteYPositionReg_95 = _RAND_230[9:0];
  _RAND_231 = {1{`RANDOM}};
  spriteYPositionReg_96 = _RAND_231[9:0];
  _RAND_232 = {1{`RANDOM}};
  spriteYPositionReg_97 = _RAND_232[9:0];
  _RAND_233 = {1{`RANDOM}};
  spriteYPositionReg_98 = _RAND_233[9:0];
  _RAND_234 = {1{`RANDOM}};
  spriteYPositionReg_99 = _RAND_234[9:0];
  _RAND_235 = {1{`RANDOM}};
  spriteYPositionReg_100 = _RAND_235[9:0];
  _RAND_236 = {1{`RANDOM}};
  spriteYPositionReg_101 = _RAND_236[9:0];
  _RAND_237 = {1{`RANDOM}};
  spriteYPositionReg_102 = _RAND_237[9:0];
  _RAND_238 = {1{`RANDOM}};
  spriteYPositionReg_103 = _RAND_238[9:0];
  _RAND_239 = {1{`RANDOM}};
  spriteYPositionReg_104 = _RAND_239[9:0];
  _RAND_240 = {1{`RANDOM}};
  spriteYPositionReg_105 = _RAND_240[9:0];
  _RAND_241 = {1{`RANDOM}};
  spriteYPositionReg_106 = _RAND_241[9:0];
  _RAND_242 = {1{`RANDOM}};
  spriteYPositionReg_107 = _RAND_242[9:0];
  _RAND_243 = {1{`RANDOM}};
  spriteYPositionReg_108 = _RAND_243[9:0];
  _RAND_244 = {1{`RANDOM}};
  spriteYPositionReg_109 = _RAND_244[9:0];
  _RAND_245 = {1{`RANDOM}};
  spriteYPositionReg_110 = _RAND_245[9:0];
  _RAND_246 = {1{`RANDOM}};
  spriteYPositionReg_111 = _RAND_246[9:0];
  _RAND_247 = {1{`RANDOM}};
  spriteYPositionReg_112 = _RAND_247[9:0];
  _RAND_248 = {1{`RANDOM}};
  spriteYPositionReg_113 = _RAND_248[9:0];
  _RAND_249 = {1{`RANDOM}};
  spriteYPositionReg_114 = _RAND_249[9:0];
  _RAND_250 = {1{`RANDOM}};
  spriteYPositionReg_115 = _RAND_250[9:0];
  _RAND_251 = {1{`RANDOM}};
  spriteYPositionReg_116 = _RAND_251[9:0];
  _RAND_252 = {1{`RANDOM}};
  spriteYPositionReg_117 = _RAND_252[9:0];
  _RAND_253 = {1{`RANDOM}};
  spriteYPositionReg_118 = _RAND_253[9:0];
  _RAND_254 = {1{`RANDOM}};
  spriteYPositionReg_119 = _RAND_254[9:0];
  _RAND_255 = {1{`RANDOM}};
  spriteYPositionReg_120 = _RAND_255[9:0];
  _RAND_256 = {1{`RANDOM}};
  spriteYPositionReg_121 = _RAND_256[9:0];
  _RAND_257 = {1{`RANDOM}};
  spriteYPositionReg_122 = _RAND_257[9:0];
  _RAND_258 = {1{`RANDOM}};
  spriteYPositionReg_123 = _RAND_258[9:0];
  _RAND_259 = {1{`RANDOM}};
  spriteYPositionReg_124 = _RAND_259[9:0];
  _RAND_260 = {1{`RANDOM}};
  spriteYPositionReg_125 = _RAND_260[9:0];
  _RAND_261 = {1{`RANDOM}};
  spriteYPositionReg_126 = _RAND_261[9:0];
  _RAND_262 = {1{`RANDOM}};
  spriteYPositionReg_127 = _RAND_262[9:0];
  _RAND_263 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  spriteVisibleReg_32 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  spriteVisibleReg_33 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  spriteVisibleReg_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  spriteVisibleReg_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  spriteVisibleReg_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  spriteVisibleReg_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  spriteVisibleReg_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  spriteVisibleReg_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  spriteVisibleReg_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  spriteVisibleReg_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  spriteVisibleReg_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  spriteVisibleReg_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  spriteVisibleReg_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  spriteVisibleReg_55 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  spriteVisibleReg_56 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  spriteVisibleReg_57 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  spriteVisibleReg_61 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  spriteVisibleReg_62 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  spriteVisibleReg_63 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  spriteVisibleReg_64 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  spriteVisibleReg_65 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  spriteVisibleReg_66 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  spriteVisibleReg_70 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  spriteVisibleReg_71 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  spriteVisibleReg_72 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  spriteFlipVerticalReg_122 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  spriteFlipVerticalReg_123 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  spriteFlipVerticalReg_124 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  spriteFlipVerticalReg_125 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  spriteFlipVerticalReg_126 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  spriteFlipVerticalReg_127 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  viewBoxXReg_0 = _RAND_326[9:0];
  _RAND_327 = {1{`RANDOM}};
  missingFrameErrorReg = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  backBufferWriteErrorReg = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  viewBoxOutOfRangeErrorReg = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  newFrameStikyReg = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  _T_47 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  backTileMemoryDataRead_0_0 = _RAND_332[6:0];
  _RAND_333 = {1{`RANDOM}};
  backTileMemoryDataRead_0_1 = _RAND_333[6:0];
  _RAND_334 = {1{`RANDOM}};
  backTileMemoryDataRead_0_2 = _RAND_334[6:0];
  _RAND_335 = {1{`RANDOM}};
  backTileMemoryDataRead_0_3 = _RAND_335[6:0];
  _RAND_336 = {1{`RANDOM}};
  backTileMemoryDataRead_0_4 = _RAND_336[6:0];
  _RAND_337 = {1{`RANDOM}};
  backTileMemoryDataRead_0_5 = _RAND_337[6:0];
  _RAND_338 = {1{`RANDOM}};
  backTileMemoryDataRead_0_6 = _RAND_338[6:0];
  _RAND_339 = {1{`RANDOM}};
  backTileMemoryDataRead_0_7 = _RAND_339[6:0];
  _RAND_340 = {1{`RANDOM}};
  backTileMemoryDataRead_0_8 = _RAND_340[6:0];
  _RAND_341 = {1{`RANDOM}};
  backTileMemoryDataRead_0_9 = _RAND_341[6:0];
  _RAND_342 = {1{`RANDOM}};
  backTileMemoryDataRead_0_10 = _RAND_342[6:0];
  _RAND_343 = {1{`RANDOM}};
  backTileMemoryDataRead_0_11 = _RAND_343[6:0];
  _RAND_344 = {1{`RANDOM}};
  backTileMemoryDataRead_0_12 = _RAND_344[6:0];
  _RAND_345 = {1{`RANDOM}};
  backTileMemoryDataRead_0_13 = _RAND_345[6:0];
  _RAND_346 = {1{`RANDOM}};
  backTileMemoryDataRead_0_14 = _RAND_346[6:0];
  _RAND_347 = {1{`RANDOM}};
  backTileMemoryDataRead_0_15 = _RAND_347[6:0];
  _RAND_348 = {1{`RANDOM}};
  backTileMemoryDataRead_0_16 = _RAND_348[6:0];
  _RAND_349 = {1{`RANDOM}};
  backTileMemoryDataRead_0_17 = _RAND_349[6:0];
  _RAND_350 = {1{`RANDOM}};
  backTileMemoryDataRead_0_18 = _RAND_350[6:0];
  _RAND_351 = {1{`RANDOM}};
  backTileMemoryDataRead_0_19 = _RAND_351[6:0];
  _RAND_352 = {1{`RANDOM}};
  backTileMemoryDataRead_0_20 = _RAND_352[6:0];
  _RAND_353 = {1{`RANDOM}};
  backTileMemoryDataRead_0_21 = _RAND_353[6:0];
  _RAND_354 = {1{`RANDOM}};
  backTileMemoryDataRead_0_22 = _RAND_354[6:0];
  _RAND_355 = {1{`RANDOM}};
  backTileMemoryDataRead_0_23 = _RAND_355[6:0];
  _RAND_356 = {1{`RANDOM}};
  backTileMemoryDataRead_0_24 = _RAND_356[6:0];
  _RAND_357 = {1{`RANDOM}};
  backTileMemoryDataRead_0_25 = _RAND_357[6:0];
  _RAND_358 = {1{`RANDOM}};
  backTileMemoryDataRead_0_26 = _RAND_358[6:0];
  _RAND_359 = {1{`RANDOM}};
  backTileMemoryDataRead_0_27 = _RAND_359[6:0];
  _RAND_360 = {1{`RANDOM}};
  backTileMemoryDataRead_0_28 = _RAND_360[6:0];
  _RAND_361 = {1{`RANDOM}};
  backTileMemoryDataRead_0_29 = _RAND_361[6:0];
  _RAND_362 = {1{`RANDOM}};
  backTileMemoryDataRead_0_30 = _RAND_362[6:0];
  _RAND_363 = {1{`RANDOM}};
  backTileMemoryDataRead_0_31 = _RAND_363[6:0];
  _RAND_364 = {1{`RANDOM}};
  backTileMemoryDataRead_1_0 = _RAND_364[6:0];
  _RAND_365 = {1{`RANDOM}};
  backTileMemoryDataRead_1_1 = _RAND_365[6:0];
  _RAND_366 = {1{`RANDOM}};
  backTileMemoryDataRead_1_2 = _RAND_366[6:0];
  _RAND_367 = {1{`RANDOM}};
  backTileMemoryDataRead_1_3 = _RAND_367[6:0];
  _RAND_368 = {1{`RANDOM}};
  backTileMemoryDataRead_1_4 = _RAND_368[6:0];
  _RAND_369 = {1{`RANDOM}};
  backTileMemoryDataRead_1_5 = _RAND_369[6:0];
  _RAND_370 = {1{`RANDOM}};
  backTileMemoryDataRead_1_6 = _RAND_370[6:0];
  _RAND_371 = {1{`RANDOM}};
  backTileMemoryDataRead_1_7 = _RAND_371[6:0];
  _RAND_372 = {1{`RANDOM}};
  backTileMemoryDataRead_1_8 = _RAND_372[6:0];
  _RAND_373 = {1{`RANDOM}};
  backTileMemoryDataRead_1_9 = _RAND_373[6:0];
  _RAND_374 = {1{`RANDOM}};
  backTileMemoryDataRead_1_10 = _RAND_374[6:0];
  _RAND_375 = {1{`RANDOM}};
  backTileMemoryDataRead_1_11 = _RAND_375[6:0];
  _RAND_376 = {1{`RANDOM}};
  backTileMemoryDataRead_1_12 = _RAND_376[6:0];
  _RAND_377 = {1{`RANDOM}};
  backTileMemoryDataRead_1_13 = _RAND_377[6:0];
  _RAND_378 = {1{`RANDOM}};
  backTileMemoryDataRead_1_14 = _RAND_378[6:0];
  _RAND_379 = {1{`RANDOM}};
  backTileMemoryDataRead_1_15 = _RAND_379[6:0];
  _RAND_380 = {1{`RANDOM}};
  backTileMemoryDataRead_1_16 = _RAND_380[6:0];
  _RAND_381 = {1{`RANDOM}};
  backTileMemoryDataRead_1_17 = _RAND_381[6:0];
  _RAND_382 = {1{`RANDOM}};
  backTileMemoryDataRead_1_18 = _RAND_382[6:0];
  _RAND_383 = {1{`RANDOM}};
  backTileMemoryDataRead_1_19 = _RAND_383[6:0];
  _RAND_384 = {1{`RANDOM}};
  backTileMemoryDataRead_1_20 = _RAND_384[6:0];
  _RAND_385 = {1{`RANDOM}};
  backTileMemoryDataRead_1_21 = _RAND_385[6:0];
  _RAND_386 = {1{`RANDOM}};
  backTileMemoryDataRead_1_22 = _RAND_386[6:0];
  _RAND_387 = {1{`RANDOM}};
  backTileMemoryDataRead_1_23 = _RAND_387[6:0];
  _RAND_388 = {1{`RANDOM}};
  backTileMemoryDataRead_1_24 = _RAND_388[6:0];
  _RAND_389 = {1{`RANDOM}};
  backTileMemoryDataRead_1_25 = _RAND_389[6:0];
  _RAND_390 = {1{`RANDOM}};
  backTileMemoryDataRead_1_26 = _RAND_390[6:0];
  _RAND_391 = {1{`RANDOM}};
  backTileMemoryDataRead_1_27 = _RAND_391[6:0];
  _RAND_392 = {1{`RANDOM}};
  backTileMemoryDataRead_1_28 = _RAND_392[6:0];
  _RAND_393 = {1{`RANDOM}};
  backTileMemoryDataRead_1_29 = _RAND_393[6:0];
  _RAND_394 = {1{`RANDOM}};
  backTileMemoryDataRead_1_30 = _RAND_394[6:0];
  _RAND_395 = {1{`RANDOM}};
  backTileMemoryDataRead_1_31 = _RAND_395[6:0];
  _RAND_396 = {1{`RANDOM}};
  backMemoryCopyCounter = _RAND_396[11:0];
  _RAND_397 = {1{`RANDOM}};
  copyEnabledReg = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  _T_377 = _RAND_398[10:0];
  _RAND_399 = {1{`RANDOM}};
  _T_379 = _RAND_399[10:0];
  _RAND_400 = {1{`RANDOM}};
  _T_382 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  _T_383 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  _T_386 = _RAND_402[4:0];
  _RAND_403 = {1{`RANDOM}};
  _T_389 = _RAND_403[10:0];
  _RAND_404 = {1{`RANDOM}};
  _T_397 = _RAND_404[10:0];
  _RAND_405 = {1{`RANDOM}};
  _T_399 = _RAND_405[10:0];
  _RAND_406 = {1{`RANDOM}};
  _T_402 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  _T_403 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  _T_406 = _RAND_408[4:0];
  _RAND_409 = {1{`RANDOM}};
  _T_409 = _RAND_409[10:0];
  _RAND_410 = {1{`RANDOM}};
  _T_416 = _RAND_410[4:0];
  _RAND_411 = {1{`RANDOM}};
  _T_419 = _RAND_411[4:0];
  _RAND_412 = {1{`RANDOM}};
  pixelColorBack = _RAND_412[5:0];
  _RAND_413 = {1{`RANDOM}};
  inSpriteX_0 = _RAND_413[11:0];
  _RAND_414 = {1{`RANDOM}};
  _T_444 = _RAND_414[11:0];
  _RAND_415 = {1{`RANDOM}};
  inSpriteX_1 = _RAND_415[11:0];
  _RAND_416 = {1{`RANDOM}};
  _T_563 = _RAND_416[11:0];
  _RAND_417 = {1{`RANDOM}};
  inSpriteX_2 = _RAND_417[11:0];
  _RAND_418 = {1{`RANDOM}};
  _T_682 = _RAND_418[11:0];
  _RAND_419 = {1{`RANDOM}};
  inSpriteX_3 = _RAND_419[11:0];
  _RAND_420 = {1{`RANDOM}};
  _T_801 = _RAND_420[11:0];
  _RAND_421 = {1{`RANDOM}};
  inSpriteX_4 = _RAND_421[11:0];
  _RAND_422 = {1{`RANDOM}};
  _T_920 = _RAND_422[11:0];
  _RAND_423 = {1{`RANDOM}};
  inSpriteX_5 = _RAND_423[11:0];
  _RAND_424 = {1{`RANDOM}};
  _T_1039 = _RAND_424[11:0];
  _RAND_425 = {1{`RANDOM}};
  inSpriteX_6 = _RAND_425[11:0];
  _RAND_426 = {1{`RANDOM}};
  _T_1158 = _RAND_426[11:0];
  _RAND_427 = {1{`RANDOM}};
  inSpriteX_7 = _RAND_427[11:0];
  _RAND_428 = {1{`RANDOM}};
  _T_1277 = _RAND_428[11:0];
  _RAND_429 = {1{`RANDOM}};
  inSpriteX_8 = _RAND_429[11:0];
  _RAND_430 = {1{`RANDOM}};
  _T_1396 = _RAND_430[11:0];
  _RAND_431 = {1{`RANDOM}};
  inSpriteX_9 = _RAND_431[11:0];
  _RAND_432 = {1{`RANDOM}};
  _T_1515 = _RAND_432[11:0];
  _RAND_433 = {1{`RANDOM}};
  inSpriteX_10 = _RAND_433[11:0];
  _RAND_434 = {1{`RANDOM}};
  _T_1634 = _RAND_434[11:0];
  _RAND_435 = {1{`RANDOM}};
  inSpriteX_11 = _RAND_435[11:0];
  _RAND_436 = {1{`RANDOM}};
  _T_1753 = _RAND_436[11:0];
  _RAND_437 = {1{`RANDOM}};
  inSpriteX_12 = _RAND_437[11:0];
  _RAND_438 = {1{`RANDOM}};
  _T_1872 = _RAND_438[11:0];
  _RAND_439 = {1{`RANDOM}};
  inSpriteX_13 = _RAND_439[11:0];
  _RAND_440 = {1{`RANDOM}};
  _T_1991 = _RAND_440[11:0];
  _RAND_441 = {1{`RANDOM}};
  inSpriteX_14 = _RAND_441[11:0];
  _RAND_442 = {1{`RANDOM}};
  _T_2110 = _RAND_442[11:0];
  _RAND_443 = {1{`RANDOM}};
  inSpriteX_15 = _RAND_443[11:0];
  _RAND_444 = {1{`RANDOM}};
  _T_2229 = _RAND_444[11:0];
  _RAND_445 = {1{`RANDOM}};
  inSpriteX_16 = _RAND_445[11:0];
  _RAND_446 = {1{`RANDOM}};
  _T_2348 = _RAND_446[11:0];
  _RAND_447 = {1{`RANDOM}};
  inSpriteX_17 = _RAND_447[11:0];
  _RAND_448 = {1{`RANDOM}};
  _T_2467 = _RAND_448[11:0];
  _RAND_449 = {1{`RANDOM}};
  inSpriteX_18 = _RAND_449[11:0];
  _RAND_450 = {1{`RANDOM}};
  _T_2586 = _RAND_450[11:0];
  _RAND_451 = {1{`RANDOM}};
  inSpriteX_19 = _RAND_451[11:0];
  _RAND_452 = {1{`RANDOM}};
  _T_2705 = _RAND_452[11:0];
  _RAND_453 = {1{`RANDOM}};
  inSpriteX_20 = _RAND_453[11:0];
  _RAND_454 = {1{`RANDOM}};
  _T_2824 = _RAND_454[11:0];
  _RAND_455 = {1{`RANDOM}};
  inSpriteX_21 = _RAND_455[11:0];
  _RAND_456 = {1{`RANDOM}};
  _T_2943 = _RAND_456[11:0];
  _RAND_457 = {1{`RANDOM}};
  inSpriteX_22 = _RAND_457[11:0];
  _RAND_458 = {1{`RANDOM}};
  _T_3062 = _RAND_458[11:0];
  _RAND_459 = {1{`RANDOM}};
  inSpriteX_23 = _RAND_459[11:0];
  _RAND_460 = {1{`RANDOM}};
  _T_3181 = _RAND_460[11:0];
  _RAND_461 = {1{`RANDOM}};
  inSpriteX_24 = _RAND_461[11:0];
  _RAND_462 = {1{`RANDOM}};
  _T_3300 = _RAND_462[11:0];
  _RAND_463 = {1{`RANDOM}};
  inSpriteX_25 = _RAND_463[11:0];
  _RAND_464 = {1{`RANDOM}};
  _T_3419 = _RAND_464[11:0];
  _RAND_465 = {1{`RANDOM}};
  inSpriteX_26 = _RAND_465[11:0];
  _RAND_466 = {1{`RANDOM}};
  _T_3538 = _RAND_466[11:0];
  _RAND_467 = {1{`RANDOM}};
  inSpriteX_27 = _RAND_467[11:0];
  _RAND_468 = {1{`RANDOM}};
  _T_3657 = _RAND_468[11:0];
  _RAND_469 = {1{`RANDOM}};
  inSpriteX_28 = _RAND_469[11:0];
  _RAND_470 = {1{`RANDOM}};
  _T_3776 = _RAND_470[11:0];
  _RAND_471 = {1{`RANDOM}};
  inSpriteX_29 = _RAND_471[11:0];
  _RAND_472 = {1{`RANDOM}};
  _T_3895 = _RAND_472[11:0];
  _RAND_473 = {1{`RANDOM}};
  inSpriteX_30 = _RAND_473[11:0];
  _RAND_474 = {1{`RANDOM}};
  _T_4014 = _RAND_474[11:0];
  _RAND_475 = {1{`RANDOM}};
  inSpriteX_31 = _RAND_475[11:0];
  _RAND_476 = {1{`RANDOM}};
  _T_4133 = _RAND_476[11:0];
  _RAND_477 = {1{`RANDOM}};
  inSpriteX_32 = _RAND_477[11:0];
  _RAND_478 = {1{`RANDOM}};
  _T_4252 = _RAND_478[11:0];
  _RAND_479 = {1{`RANDOM}};
  inSpriteX_33 = _RAND_479[11:0];
  _RAND_480 = {1{`RANDOM}};
  _T_4371 = _RAND_480[11:0];
  _RAND_481 = {1{`RANDOM}};
  inSpriteX_34 = _RAND_481[11:0];
  _RAND_482 = {1{`RANDOM}};
  _T_4490 = _RAND_482[11:0];
  _RAND_483 = {1{`RANDOM}};
  inSpriteX_35 = _RAND_483[11:0];
  _RAND_484 = {1{`RANDOM}};
  _T_4609 = _RAND_484[11:0];
  _RAND_485 = {1{`RANDOM}};
  inSpriteX_36 = _RAND_485[11:0];
  _RAND_486 = {1{`RANDOM}};
  _T_4728 = _RAND_486[11:0];
  _RAND_487 = {1{`RANDOM}};
  inSpriteX_37 = _RAND_487[11:0];
  _RAND_488 = {1{`RANDOM}};
  _T_4847 = _RAND_488[11:0];
  _RAND_489 = {1{`RANDOM}};
  inSpriteX_38 = _RAND_489[11:0];
  _RAND_490 = {1{`RANDOM}};
  _T_4966 = _RAND_490[11:0];
  _RAND_491 = {1{`RANDOM}};
  inSpriteX_39 = _RAND_491[11:0];
  _RAND_492 = {1{`RANDOM}};
  _T_5085 = _RAND_492[11:0];
  _RAND_493 = {1{`RANDOM}};
  inSpriteX_40 = _RAND_493[11:0];
  _RAND_494 = {1{`RANDOM}};
  _T_5204 = _RAND_494[11:0];
  _RAND_495 = {1{`RANDOM}};
  inSpriteX_41 = _RAND_495[11:0];
  _RAND_496 = {1{`RANDOM}};
  _T_5323 = _RAND_496[11:0];
  _RAND_497 = {1{`RANDOM}};
  inSpriteX_42 = _RAND_497[11:0];
  _RAND_498 = {1{`RANDOM}};
  _T_5442 = _RAND_498[11:0];
  _RAND_499 = {1{`RANDOM}};
  inSpriteX_43 = _RAND_499[11:0];
  _RAND_500 = {1{`RANDOM}};
  _T_5561 = _RAND_500[11:0];
  _RAND_501 = {1{`RANDOM}};
  inSpriteX_44 = _RAND_501[11:0];
  _RAND_502 = {1{`RANDOM}};
  _T_5680 = _RAND_502[11:0];
  _RAND_503 = {1{`RANDOM}};
  inSpriteX_45 = _RAND_503[11:0];
  _RAND_504 = {1{`RANDOM}};
  _T_5799 = _RAND_504[11:0];
  _RAND_505 = {1{`RANDOM}};
  inSpriteX_46 = _RAND_505[11:0];
  _RAND_506 = {1{`RANDOM}};
  _T_5918 = _RAND_506[11:0];
  _RAND_507 = {1{`RANDOM}};
  inSpriteX_47 = _RAND_507[11:0];
  _RAND_508 = {1{`RANDOM}};
  _T_6037 = _RAND_508[11:0];
  _RAND_509 = {1{`RANDOM}};
  inSpriteX_48 = _RAND_509[11:0];
  _RAND_510 = {1{`RANDOM}};
  _T_6156 = _RAND_510[11:0];
  _RAND_511 = {1{`RANDOM}};
  inSpriteX_49 = _RAND_511[11:0];
  _RAND_512 = {1{`RANDOM}};
  _T_6275 = _RAND_512[11:0];
  _RAND_513 = {1{`RANDOM}};
  inSpriteX_50 = _RAND_513[11:0];
  _RAND_514 = {1{`RANDOM}};
  _T_6394 = _RAND_514[11:0];
  _RAND_515 = {1{`RANDOM}};
  inSpriteX_51 = _RAND_515[11:0];
  _RAND_516 = {1{`RANDOM}};
  _T_6513 = _RAND_516[11:0];
  _RAND_517 = {1{`RANDOM}};
  inSpriteX_52 = _RAND_517[11:0];
  _RAND_518 = {1{`RANDOM}};
  _T_6632 = _RAND_518[11:0];
  _RAND_519 = {1{`RANDOM}};
  inSpriteX_53 = _RAND_519[11:0];
  _RAND_520 = {1{`RANDOM}};
  _T_6751 = _RAND_520[11:0];
  _RAND_521 = {1{`RANDOM}};
  inSpriteX_54 = _RAND_521[11:0];
  _RAND_522 = {1{`RANDOM}};
  _T_6870 = _RAND_522[11:0];
  _RAND_523 = {1{`RANDOM}};
  inSpriteX_55 = _RAND_523[11:0];
  _RAND_524 = {1{`RANDOM}};
  _T_6989 = _RAND_524[11:0];
  _RAND_525 = {1{`RANDOM}};
  inSpriteX_56 = _RAND_525[11:0];
  _RAND_526 = {1{`RANDOM}};
  _T_7108 = _RAND_526[11:0];
  _RAND_527 = {1{`RANDOM}};
  inSpriteX_57 = _RAND_527[11:0];
  _RAND_528 = {1{`RANDOM}};
  _T_7227 = _RAND_528[11:0];
  _RAND_529 = {1{`RANDOM}};
  inSpriteX_58 = _RAND_529[11:0];
  _RAND_530 = {1{`RANDOM}};
  _T_7346 = _RAND_530[11:0];
  _RAND_531 = {1{`RANDOM}};
  inSpriteX_59 = _RAND_531[11:0];
  _RAND_532 = {1{`RANDOM}};
  _T_7465 = _RAND_532[11:0];
  _RAND_533 = {1{`RANDOM}};
  inSpriteX_60 = _RAND_533[11:0];
  _RAND_534 = {1{`RANDOM}};
  _T_7584 = _RAND_534[11:0];
  _RAND_535 = {1{`RANDOM}};
  inSpriteX_61 = _RAND_535[11:0];
  _RAND_536 = {1{`RANDOM}};
  _T_7703 = _RAND_536[11:0];
  _RAND_537 = {1{`RANDOM}};
  inSpriteX_62 = _RAND_537[11:0];
  _RAND_538 = {1{`RANDOM}};
  _T_7822 = _RAND_538[11:0];
  _RAND_539 = {1{`RANDOM}};
  inSpriteX_63 = _RAND_539[11:0];
  _RAND_540 = {1{`RANDOM}};
  _T_7941 = _RAND_540[11:0];
  _RAND_541 = {1{`RANDOM}};
  inSpriteX_64 = _RAND_541[11:0];
  _RAND_542 = {1{`RANDOM}};
  _T_8060 = _RAND_542[11:0];
  _RAND_543 = {1{`RANDOM}};
  inSpriteX_65 = _RAND_543[11:0];
  _RAND_544 = {1{`RANDOM}};
  _T_8179 = _RAND_544[11:0];
  _RAND_545 = {1{`RANDOM}};
  inSpriteX_66 = _RAND_545[11:0];
  _RAND_546 = {1{`RANDOM}};
  _T_8298 = _RAND_546[11:0];
  _RAND_547 = {1{`RANDOM}};
  inSpriteX_67 = _RAND_547[11:0];
  _RAND_548 = {1{`RANDOM}};
  _T_8417 = _RAND_548[11:0];
  _RAND_549 = {1{`RANDOM}};
  inSpriteX_68 = _RAND_549[11:0];
  _RAND_550 = {1{`RANDOM}};
  _T_8536 = _RAND_550[11:0];
  _RAND_551 = {1{`RANDOM}};
  inSpriteX_69 = _RAND_551[11:0];
  _RAND_552 = {1{`RANDOM}};
  _T_8655 = _RAND_552[11:0];
  _RAND_553 = {1{`RANDOM}};
  inSpriteX_70 = _RAND_553[11:0];
  _RAND_554 = {1{`RANDOM}};
  _T_8774 = _RAND_554[11:0];
  _RAND_555 = {1{`RANDOM}};
  inSpriteX_71 = _RAND_555[11:0];
  _RAND_556 = {1{`RANDOM}};
  _T_8893 = _RAND_556[11:0];
  _RAND_557 = {1{`RANDOM}};
  inSpriteX_72 = _RAND_557[11:0];
  _RAND_558 = {1{`RANDOM}};
  _T_9012 = _RAND_558[11:0];
  _RAND_559 = {1{`RANDOM}};
  inSpriteX_73 = _RAND_559[11:0];
  _RAND_560 = {1{`RANDOM}};
  _T_9131 = _RAND_560[11:0];
  _RAND_561 = {1{`RANDOM}};
  inSpriteX_74 = _RAND_561[11:0];
  _RAND_562 = {1{`RANDOM}};
  _T_9250 = _RAND_562[11:0];
  _RAND_563 = {1{`RANDOM}};
  inSpriteX_75 = _RAND_563[11:0];
  _RAND_564 = {1{`RANDOM}};
  _T_9369 = _RAND_564[11:0];
  _RAND_565 = {1{`RANDOM}};
  inSpriteX_76 = _RAND_565[11:0];
  _RAND_566 = {1{`RANDOM}};
  _T_9488 = _RAND_566[11:0];
  _RAND_567 = {1{`RANDOM}};
  inSpriteX_77 = _RAND_567[11:0];
  _RAND_568 = {1{`RANDOM}};
  _T_9607 = _RAND_568[11:0];
  _RAND_569 = {1{`RANDOM}};
  inSpriteX_78 = _RAND_569[11:0];
  _RAND_570 = {1{`RANDOM}};
  _T_9726 = _RAND_570[11:0];
  _RAND_571 = {1{`RANDOM}};
  inSpriteX_79 = _RAND_571[11:0];
  _RAND_572 = {1{`RANDOM}};
  _T_9845 = _RAND_572[11:0];
  _RAND_573 = {1{`RANDOM}};
  inSpriteX_80 = _RAND_573[11:0];
  _RAND_574 = {1{`RANDOM}};
  _T_9964 = _RAND_574[11:0];
  _RAND_575 = {1{`RANDOM}};
  inSpriteX_81 = _RAND_575[11:0];
  _RAND_576 = {1{`RANDOM}};
  _T_10083 = _RAND_576[11:0];
  _RAND_577 = {1{`RANDOM}};
  inSpriteX_82 = _RAND_577[11:0];
  _RAND_578 = {1{`RANDOM}};
  _T_10202 = _RAND_578[11:0];
  _RAND_579 = {1{`RANDOM}};
  inSpriteX_83 = _RAND_579[11:0];
  _RAND_580 = {1{`RANDOM}};
  _T_10321 = _RAND_580[11:0];
  _RAND_581 = {1{`RANDOM}};
  inSpriteX_84 = _RAND_581[11:0];
  _RAND_582 = {1{`RANDOM}};
  _T_10440 = _RAND_582[11:0];
  _RAND_583 = {1{`RANDOM}};
  inSpriteX_85 = _RAND_583[11:0];
  _RAND_584 = {1{`RANDOM}};
  _T_10559 = _RAND_584[11:0];
  _RAND_585 = {1{`RANDOM}};
  inSpriteX_86 = _RAND_585[11:0];
  _RAND_586 = {1{`RANDOM}};
  _T_10678 = _RAND_586[11:0];
  _RAND_587 = {1{`RANDOM}};
  inSpriteX_87 = _RAND_587[11:0];
  _RAND_588 = {1{`RANDOM}};
  _T_10797 = _RAND_588[11:0];
  _RAND_589 = {1{`RANDOM}};
  inSpriteX_88 = _RAND_589[11:0];
  _RAND_590 = {1{`RANDOM}};
  _T_10916 = _RAND_590[11:0];
  _RAND_591 = {1{`RANDOM}};
  inSpriteX_89 = _RAND_591[11:0];
  _RAND_592 = {1{`RANDOM}};
  _T_11035 = _RAND_592[11:0];
  _RAND_593 = {1{`RANDOM}};
  inSpriteX_90 = _RAND_593[11:0];
  _RAND_594 = {1{`RANDOM}};
  _T_11154 = _RAND_594[11:0];
  _RAND_595 = {1{`RANDOM}};
  inSpriteX_91 = _RAND_595[11:0];
  _RAND_596 = {1{`RANDOM}};
  _T_11273 = _RAND_596[11:0];
  _RAND_597 = {1{`RANDOM}};
  inSpriteX_92 = _RAND_597[11:0];
  _RAND_598 = {1{`RANDOM}};
  _T_11392 = _RAND_598[11:0];
  _RAND_599 = {1{`RANDOM}};
  inSpriteX_93 = _RAND_599[11:0];
  _RAND_600 = {1{`RANDOM}};
  _T_11511 = _RAND_600[11:0];
  _RAND_601 = {1{`RANDOM}};
  inSpriteX_94 = _RAND_601[11:0];
  _RAND_602 = {1{`RANDOM}};
  _T_11630 = _RAND_602[11:0];
  _RAND_603 = {1{`RANDOM}};
  inSpriteX_95 = _RAND_603[11:0];
  _RAND_604 = {1{`RANDOM}};
  _T_11749 = _RAND_604[11:0];
  _RAND_605 = {1{`RANDOM}};
  inSpriteX_96 = _RAND_605[11:0];
  _RAND_606 = {1{`RANDOM}};
  _T_11868 = _RAND_606[11:0];
  _RAND_607 = {1{`RANDOM}};
  inSpriteX_97 = _RAND_607[11:0];
  _RAND_608 = {1{`RANDOM}};
  _T_11987 = _RAND_608[11:0];
  _RAND_609 = {1{`RANDOM}};
  inSpriteX_98 = _RAND_609[11:0];
  _RAND_610 = {1{`RANDOM}};
  _T_12106 = _RAND_610[11:0];
  _RAND_611 = {1{`RANDOM}};
  inSpriteX_99 = _RAND_611[11:0];
  _RAND_612 = {1{`RANDOM}};
  _T_12225 = _RAND_612[11:0];
  _RAND_613 = {1{`RANDOM}};
  inSpriteX_100 = _RAND_613[11:0];
  _RAND_614 = {1{`RANDOM}};
  _T_12344 = _RAND_614[11:0];
  _RAND_615 = {1{`RANDOM}};
  inSpriteX_101 = _RAND_615[11:0];
  _RAND_616 = {1{`RANDOM}};
  _T_12463 = _RAND_616[11:0];
  _RAND_617 = {1{`RANDOM}};
  inSpriteX_102 = _RAND_617[11:0];
  _RAND_618 = {1{`RANDOM}};
  _T_12582 = _RAND_618[11:0];
  _RAND_619 = {1{`RANDOM}};
  inSpriteX_103 = _RAND_619[11:0];
  _RAND_620 = {1{`RANDOM}};
  _T_12701 = _RAND_620[11:0];
  _RAND_621 = {1{`RANDOM}};
  inSpriteX_104 = _RAND_621[11:0];
  _RAND_622 = {1{`RANDOM}};
  _T_12820 = _RAND_622[11:0];
  _RAND_623 = {1{`RANDOM}};
  inSpriteX_105 = _RAND_623[11:0];
  _RAND_624 = {1{`RANDOM}};
  _T_12939 = _RAND_624[11:0];
  _RAND_625 = {1{`RANDOM}};
  inSpriteX_106 = _RAND_625[11:0];
  _RAND_626 = {1{`RANDOM}};
  _T_13058 = _RAND_626[11:0];
  _RAND_627 = {1{`RANDOM}};
  inSpriteX_107 = _RAND_627[11:0];
  _RAND_628 = {1{`RANDOM}};
  _T_13177 = _RAND_628[11:0];
  _RAND_629 = {1{`RANDOM}};
  inSpriteX_108 = _RAND_629[11:0];
  _RAND_630 = {1{`RANDOM}};
  _T_13296 = _RAND_630[11:0];
  _RAND_631 = {1{`RANDOM}};
  inSpriteX_109 = _RAND_631[11:0];
  _RAND_632 = {1{`RANDOM}};
  _T_13415 = _RAND_632[11:0];
  _RAND_633 = {1{`RANDOM}};
  inSpriteX_110 = _RAND_633[11:0];
  _RAND_634 = {1{`RANDOM}};
  _T_13534 = _RAND_634[11:0];
  _RAND_635 = {1{`RANDOM}};
  inSpriteX_111 = _RAND_635[11:0];
  _RAND_636 = {1{`RANDOM}};
  _T_13653 = _RAND_636[11:0];
  _RAND_637 = {1{`RANDOM}};
  inSpriteX_112 = _RAND_637[11:0];
  _RAND_638 = {1{`RANDOM}};
  _T_13772 = _RAND_638[11:0];
  _RAND_639 = {1{`RANDOM}};
  inSpriteX_113 = _RAND_639[11:0];
  _RAND_640 = {1{`RANDOM}};
  _T_13891 = _RAND_640[11:0];
  _RAND_641 = {1{`RANDOM}};
  inSpriteX_114 = _RAND_641[11:0];
  _RAND_642 = {1{`RANDOM}};
  _T_14010 = _RAND_642[11:0];
  _RAND_643 = {1{`RANDOM}};
  inSpriteX_115 = _RAND_643[11:0];
  _RAND_644 = {1{`RANDOM}};
  _T_14129 = _RAND_644[11:0];
  _RAND_645 = {1{`RANDOM}};
  inSpriteX_116 = _RAND_645[11:0];
  _RAND_646 = {1{`RANDOM}};
  _T_14248 = _RAND_646[11:0];
  _RAND_647 = {1{`RANDOM}};
  inSpriteX_117 = _RAND_647[11:0];
  _RAND_648 = {1{`RANDOM}};
  _T_14367 = _RAND_648[11:0];
  _RAND_649 = {1{`RANDOM}};
  inSpriteX_118 = _RAND_649[11:0];
  _RAND_650 = {1{`RANDOM}};
  _T_14486 = _RAND_650[11:0];
  _RAND_651 = {1{`RANDOM}};
  inSpriteX_119 = _RAND_651[11:0];
  _RAND_652 = {1{`RANDOM}};
  _T_14605 = _RAND_652[11:0];
  _RAND_653 = {1{`RANDOM}};
  inSpriteX_120 = _RAND_653[11:0];
  _RAND_654 = {1{`RANDOM}};
  _T_14724 = _RAND_654[11:0];
  _RAND_655 = {1{`RANDOM}};
  inSpriteX_121 = _RAND_655[11:0];
  _RAND_656 = {1{`RANDOM}};
  _T_14843 = _RAND_656[11:0];
  _RAND_657 = {1{`RANDOM}};
  inSpriteX_122 = _RAND_657[11:0];
  _RAND_658 = {1{`RANDOM}};
  _T_14962 = _RAND_658[11:0];
  _RAND_659 = {1{`RANDOM}};
  inSpriteX_123 = _RAND_659[11:0];
  _RAND_660 = {1{`RANDOM}};
  _T_15081 = _RAND_660[11:0];
  _RAND_661 = {1{`RANDOM}};
  inSpriteX_124 = _RAND_661[11:0];
  _RAND_662 = {1{`RANDOM}};
  _T_15200 = _RAND_662[11:0];
  _RAND_663 = {1{`RANDOM}};
  inSpriteX_125 = _RAND_663[11:0];
  _RAND_664 = {1{`RANDOM}};
  _T_15319 = _RAND_664[11:0];
  _RAND_665 = {1{`RANDOM}};
  inSpriteX_126 = _RAND_665[11:0];
  _RAND_666 = {1{`RANDOM}};
  _T_15438 = _RAND_666[11:0];
  _RAND_667 = {1{`RANDOM}};
  inSpriteX_127 = _RAND_667[11:0];
  _RAND_668 = {1{`RANDOM}};
  _T_15557 = _RAND_668[11:0];
  _RAND_669 = {1{`RANDOM}};
  _T_15660_0 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  _T_15660_1 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  _T_15660_2 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  _T_15662_0 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  _T_15662_1 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  _T_15662_2 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  _T_15664_0 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  _T_15664_1 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  _T_15664_2 = _RAND_677[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ScaleCounterReg <= 2'h0;
    end else if (run) begin
      if (_T) begin
        ScaleCounterReg <= 2'h0;
      end else begin
        ScaleCounterReg <= _T_8;
      end
    end
    if (reset) begin
      CounterXReg <= 10'h0;
    end else if (run) begin
      if (_T) begin
        if (_T_1) begin
          CounterXReg <= 10'h0;
        end else begin
          CounterXReg <= _T_6;
        end
      end
    end
    if (reset) begin
      CounterYReg <= 10'h0;
    end else if (run) begin
      if (_T) begin
        if (_T_1) begin
          if (_T_2) begin
            CounterYReg <= 10'h0;
          end else begin
            CounterYReg <= _T_4;
          end
        end
      end
    end
    if (reset) begin
      backMemoryRestoreCounter <= 12'h0;
    end else if (restoreEnabled) begin
      backMemoryRestoreCounter <= _T_374;
    end
    _T_14_0 <= _T_14_1;
    _T_14_1 <= _T_14_2;
    _T_14_2 <= _T_14_3;
    _T_14_3 <= ~Hsync;
    _T_16_0 <= _T_16_1;
    _T_16_1 <= _T_16_2;
    _T_16_2 <= _T_16_3;
    _T_16_3 <= ~Vsync;
    if (reset) begin
      frameClockCount <= 21'h0;
    end else if (_T_19) begin
      frameClockCount <= 21'h0;
    end else begin
      frameClockCount <= _T_21;
    end
    if (reset) begin
      spriteXPositionReg_0 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_0 <= io_spriteXPosition_0;
    end
    if (reset) begin
      spriteXPositionReg_1 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_1 <= io_spriteXPosition_1;
    end
    if (reset) begin
      spriteXPositionReg_2 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_2 <= io_spriteXPosition_2;
    end
    if (reset) begin
      spriteXPositionReg_3 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_3 <= io_spriteXPosition_3;
    end
    if (reset) begin
      spriteXPositionReg_4 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_4 <= io_spriteXPosition_4;
    end
    if (reset) begin
      spriteXPositionReg_5 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_5 <= io_spriteXPosition_5;
    end
    if (reset) begin
      spriteXPositionReg_6 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_6 <= io_spriteXPosition_6;
    end
    if (reset) begin
      spriteXPositionReg_7 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_7 <= io_spriteXPosition_7;
    end
    if (reset) begin
      spriteXPositionReg_8 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_8 <= io_spriteXPosition_8;
    end
    if (reset) begin
      spriteXPositionReg_9 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_9 <= io_spriteXPosition_9;
    end
    if (reset) begin
      spriteXPositionReg_10 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_10 <= io_spriteXPosition_10;
    end
    if (reset) begin
      spriteXPositionReg_11 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_11 <= io_spriteXPosition_11;
    end
    if (reset) begin
      spriteXPositionReg_12 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_12 <= io_spriteXPosition_12;
    end
    if (reset) begin
      spriteXPositionReg_13 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_13 <= io_spriteXPosition_13;
    end
    if (reset) begin
      spriteXPositionReg_14 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_14 <= io_spriteXPosition_14;
    end
    if (reset) begin
      spriteXPositionReg_15 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_15 <= io_spriteXPosition_15;
    end
    if (reset) begin
      spriteXPositionReg_16 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_16 <= io_spriteXPosition_16;
    end
    if (reset) begin
      spriteXPositionReg_17 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_17 <= io_spriteXPosition_17;
    end
    if (reset) begin
      spriteXPositionReg_18 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_18 <= io_spriteXPosition_18;
    end
    if (reset) begin
      spriteXPositionReg_19 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_19 <= io_spriteXPosition_19;
    end
    if (reset) begin
      spriteXPositionReg_20 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_20 <= io_spriteXPosition_20;
    end
    if (reset) begin
      spriteXPositionReg_21 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_21 <= io_spriteXPosition_21;
    end
    if (reset) begin
      spriteXPositionReg_22 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_22 <= io_spriteXPosition_22;
    end
    if (reset) begin
      spriteXPositionReg_23 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_23 <= io_spriteXPosition_23;
    end
    if (reset) begin
      spriteXPositionReg_24 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_24 <= io_spriteXPosition_24;
    end
    if (reset) begin
      spriteXPositionReg_25 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_25 <= io_spriteXPosition_25;
    end
    if (reset) begin
      spriteXPositionReg_26 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_26 <= io_spriteXPosition_26;
    end
    if (reset) begin
      spriteXPositionReg_27 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_27 <= io_spriteXPosition_27;
    end
    if (reset) begin
      spriteXPositionReg_28 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_28 <= io_spriteXPosition_28;
    end
    if (reset) begin
      spriteXPositionReg_29 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_29 <= io_spriteXPosition_29;
    end
    if (reset) begin
      spriteXPositionReg_30 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_30 <= io_spriteXPosition_30;
    end
    if (reset) begin
      spriteXPositionReg_31 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_31 <= io_spriteXPosition_31;
    end
    if (reset) begin
      spriteXPositionReg_32 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_32 <= io_spriteXPosition_32;
    end
    if (reset) begin
      spriteXPositionReg_33 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_33 <= io_spriteXPosition_33;
    end
    if (reset) begin
      spriteXPositionReg_34 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_34 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_35 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_35 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_36 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_36 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_37 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_37 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_38 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_38 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_39 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_39 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_40 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_40 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_41 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_41 <= io_spriteXPosition_41;
    end
    if (reset) begin
      spriteXPositionReg_42 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_42 <= io_spriteXPosition_42;
    end
    if (reset) begin
      spriteXPositionReg_43 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_43 <= io_spriteXPosition_43;
    end
    if (reset) begin
      spriteXPositionReg_44 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_44 <= io_spriteXPosition_44;
    end
    if (reset) begin
      spriteXPositionReg_45 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_45 <= io_spriteXPosition_45;
    end
    if (reset) begin
      spriteXPositionReg_46 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_46 <= io_spriteXPosition_46;
    end
    if (reset) begin
      spriteXPositionReg_47 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_47 <= io_spriteXPosition_47;
    end
    if (reset) begin
      spriteXPositionReg_48 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_48 <= io_spriteXPosition_48;
    end
    if (reset) begin
      spriteXPositionReg_49 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_49 <= io_spriteXPosition_49;
    end
    if (reset) begin
      spriteXPositionReg_50 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_50 <= io_spriteXPosition_50;
    end
    if (reset) begin
      spriteXPositionReg_51 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_51 <= io_spriteXPosition_51;
    end
    if (reset) begin
      spriteXPositionReg_52 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_52 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_53 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_53 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_54 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_54 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_55 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_55 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_56 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_56 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_57 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_57 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_58 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_58 <= 11'sh1e0;
    end
    if (reset) begin
      spriteXPositionReg_59 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_59 <= 11'sh200;
    end
    if (reset) begin
      spriteXPositionReg_60 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_60 <= 11'sh220;
    end
    if (reset) begin
      spriteXPositionReg_61 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_61 <= 11'sh1e0;
    end
    if (reset) begin
      spriteXPositionReg_62 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_62 <= 11'sh200;
    end
    if (reset) begin
      spriteXPositionReg_63 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_63 <= 11'sh220;
    end
    if (reset) begin
      spriteXPositionReg_64 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_64 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_65 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_65 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_66 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_66 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_67 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_67 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_68 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_68 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_69 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_69 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_70 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_70 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_71 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_71 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_72 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_72 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_73 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_73 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_74 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_74 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_75 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_75 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_76 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_76 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_77 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_77 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_78 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_78 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_79 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_79 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_80 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_80 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_81 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_81 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_82 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_82 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_83 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_83 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_84 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_84 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_85 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_85 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_86 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_86 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_87 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_87 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_88 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_88 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_89 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_89 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_90 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_90 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_91 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_91 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_92 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_92 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_93 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_93 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_94 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_94 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_95 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_95 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_96 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_96 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_97 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_97 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_98 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_98 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_99 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_99 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_100 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_100 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_101 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_101 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_102 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_102 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_103 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_103 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_104 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_104 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_105 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_105 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_106 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_106 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_107 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_107 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_108 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_108 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_109 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_109 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_110 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_110 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_111 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_111 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_112 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_112 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_113 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_113 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_114 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_114 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_115 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_115 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_116 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_116 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_117 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_117 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_118 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_118 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_119 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_119 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_120 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_120 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_121 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_121 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_122 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_122 <= io_spriteXPosition_122;
    end
    if (reset) begin
      spriteXPositionReg_123 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_123 <= io_spriteXPosition_123;
    end
    if (reset) begin
      spriteXPositionReg_124 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_124 <= io_spriteXPosition_124;
    end
    if (reset) begin
      spriteXPositionReg_125 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_125 <= io_spriteXPosition_125;
    end
    if (reset) begin
      spriteXPositionReg_126 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_126 <= io_spriteXPosition_126;
    end
    if (reset) begin
      spriteXPositionReg_127 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_127 <= io_spriteXPosition_127;
    end
    if (reset) begin
      spriteYPositionReg_0 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_0 <= io_spriteYPosition_0;
    end
    if (reset) begin
      spriteYPositionReg_1 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_1 <= io_spriteYPosition_1;
    end
    if (reset) begin
      spriteYPositionReg_2 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_2 <= io_spriteYPosition_2;
    end
    if (reset) begin
      spriteYPositionReg_3 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_3 <= io_spriteYPosition_3;
    end
    if (reset) begin
      spriteYPositionReg_4 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_4 <= io_spriteYPosition_4;
    end
    if (reset) begin
      spriteYPositionReg_5 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_5 <= io_spriteYPosition_5;
    end
    if (reset) begin
      spriteYPositionReg_6 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_6 <= io_spriteYPosition_6;
    end
    if (reset) begin
      spriteYPositionReg_7 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_7 <= io_spriteYPosition_7;
    end
    if (reset) begin
      spriteYPositionReg_8 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_8 <= io_spriteYPosition_8;
    end
    if (reset) begin
      spriteYPositionReg_9 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_9 <= io_spriteYPosition_9;
    end
    if (reset) begin
      spriteYPositionReg_10 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_10 <= io_spriteYPosition_10;
    end
    if (reset) begin
      spriteYPositionReg_11 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_11 <= io_spriteYPosition_11;
    end
    if (reset) begin
      spriteYPositionReg_12 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_12 <= io_spriteYPosition_12;
    end
    if (reset) begin
      spriteYPositionReg_13 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_13 <= io_spriteYPosition_13;
    end
    if (reset) begin
      spriteYPositionReg_14 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_14 <= io_spriteYPosition_14;
    end
    if (reset) begin
      spriteYPositionReg_15 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_15 <= io_spriteYPosition_15;
    end
    if (reset) begin
      spriteYPositionReg_16 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_16 <= io_spriteYPosition_16;
    end
    if (reset) begin
      spriteYPositionReg_17 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_17 <= io_spriteYPosition_17;
    end
    if (reset) begin
      spriteYPositionReg_18 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_18 <= io_spriteYPosition_18;
    end
    if (reset) begin
      spriteYPositionReg_19 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_19 <= io_spriteYPosition_19;
    end
    if (reset) begin
      spriteYPositionReg_20 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_20 <= io_spriteYPosition_20;
    end
    if (reset) begin
      spriteYPositionReg_21 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_21 <= io_spriteYPosition_21;
    end
    if (reset) begin
      spriteYPositionReg_22 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_22 <= io_spriteYPosition_22;
    end
    if (reset) begin
      spriteYPositionReg_23 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_23 <= io_spriteYPosition_23;
    end
    if (reset) begin
      spriteYPositionReg_24 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_24 <= io_spriteYPosition_24;
    end
    if (reset) begin
      spriteYPositionReg_25 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_25 <= io_spriteYPosition_25;
    end
    if (reset) begin
      spriteYPositionReg_26 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_26 <= io_spriteYPosition_26;
    end
    if (reset) begin
      spriteYPositionReg_27 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_27 <= io_spriteYPosition_27;
    end
    if (reset) begin
      spriteYPositionReg_28 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_28 <= io_spriteYPosition_28;
    end
    if (reset) begin
      spriteYPositionReg_29 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_29 <= io_spriteYPosition_29;
    end
    if (reset) begin
      spriteYPositionReg_30 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_30 <= io_spriteYPosition_30;
    end
    if (reset) begin
      spriteYPositionReg_31 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_31 <= io_spriteYPosition_31;
    end
    if (reset) begin
      spriteYPositionReg_32 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_32 <= io_spriteYPosition_32;
    end
    if (reset) begin
      spriteYPositionReg_33 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_33 <= io_spriteYPosition_33;
    end
    if (reset) begin
      spriteYPositionReg_34 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_34 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_35 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_35 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_36 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_36 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_37 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_37 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_38 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_38 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_39 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_39 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_40 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_40 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_41 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_41 <= io_spriteYPosition_41;
    end
    if (reset) begin
      spriteYPositionReg_42 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_42 <= io_spriteYPosition_42;
    end
    if (reset) begin
      spriteYPositionReg_43 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_43 <= io_spriteYPosition_43;
    end
    if (reset) begin
      spriteYPositionReg_44 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_44 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_45 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_45 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_46 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_46 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_47 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_47 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_48 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_48 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_49 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_49 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_50 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_50 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_51 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_51 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_52 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_52 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_53 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_53 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_54 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_54 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_55 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_55 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_56 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_56 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_57 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_57 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_58 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_58 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_59 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_59 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_60 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_60 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_61 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_61 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_62 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_62 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_63 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_63 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_70 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_70 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_71 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_71 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_72 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_72 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_73 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_73 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_74 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_74 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_75 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_75 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_76 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_76 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_77 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_77 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_78 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_78 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_79 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_79 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_80 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_80 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_81 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_81 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_82 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_82 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_83 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_83 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_84 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_84 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_85 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_85 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_86 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_86 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_87 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_87 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_88 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_88 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_89 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_89 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_90 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_90 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_91 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_91 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_92 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_92 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_93 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_93 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_94 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_94 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_95 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_95 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_96 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_96 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_97 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_97 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_98 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_98 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_99 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_99 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_100 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_100 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_101 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_101 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_102 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_102 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_103 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_103 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_104 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_104 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_105 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_105 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_106 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_106 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_107 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_107 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_108 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_108 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_109 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_109 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_110 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_110 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_111 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_111 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_112 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_112 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_113 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_113 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_114 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_114 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_115 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_115 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_116 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_116 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_117 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_117 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_118 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_118 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_119 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_119 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_120 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_120 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_121 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_121 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_122 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_122 <= io_spriteYPosition_122;
    end
    if (reset) begin
      spriteYPositionReg_123 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_123 <= io_spriteYPosition_123;
    end
    if (reset) begin
      spriteYPositionReg_124 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_124 <= io_spriteYPosition_124;
    end
    if (reset) begin
      spriteYPositionReg_125 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_125 <= io_spriteYPosition_125;
    end
    if (reset) begin
      spriteYPositionReg_126 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_126 <= io_spriteYPosition_126;
    end
    if (reset) begin
      spriteYPositionReg_127 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_127 <= io_spriteYPosition_127;
    end
    spriteVisibleReg_0 <= reset | _GEN_269;
    spriteVisibleReg_1 <= reset | _GEN_270;
    spriteVisibleReg_2 <= reset | _GEN_271;
    spriteVisibleReg_3 <= reset | _GEN_272;
    spriteVisibleReg_4 <= reset | _GEN_273;
    spriteVisibleReg_5 <= reset | _GEN_274;
    spriteVisibleReg_6 <= reset | _GEN_275;
    spriteVisibleReg_7 <= reset | _GEN_276;
    spriteVisibleReg_8 <= reset | _GEN_277;
    spriteVisibleReg_9 <= reset | _GEN_278;
    spriteVisibleReg_10 <= reset | _GEN_279;
    spriteVisibleReg_11 <= reset | _GEN_280;
    spriteVisibleReg_12 <= reset | _GEN_281;
    spriteVisibleReg_13 <= reset | _GEN_282;
    spriteVisibleReg_14 <= reset | _GEN_283;
    spriteVisibleReg_15 <= reset | _GEN_284;
    spriteVisibleReg_16 <= reset | _GEN_285;
    spriteVisibleReg_17 <= reset | _GEN_286;
    spriteVisibleReg_18 <= reset | _GEN_287;
    spriteVisibleReg_19 <= reset | _GEN_288;
    spriteVisibleReg_20 <= reset | _GEN_289;
    spriteVisibleReg_21 <= reset | _GEN_290;
    spriteVisibleReg_22 <= reset | _GEN_291;
    spriteVisibleReg_23 <= reset | _GEN_292;
    spriteVisibleReg_24 <= reset | _GEN_293;
    spriteVisibleReg_25 <= reset | _GEN_294;
    spriteVisibleReg_26 <= reset | _GEN_295;
    spriteVisibleReg_27 <= reset | _GEN_296;
    spriteVisibleReg_28 <= reset | _GEN_297;
    spriteVisibleReg_29 <= reset | _GEN_298;
    spriteVisibleReg_30 <= reset | _GEN_299;
    spriteVisibleReg_31 <= reset | _GEN_300;
    spriteVisibleReg_32 <= reset | _GEN_301;
    spriteVisibleReg_33 <= reset | _GEN_302;
    spriteVisibleReg_41 <= reset | _GEN_310;
    spriteVisibleReg_42 <= reset | _GEN_311;
    spriteVisibleReg_43 <= reset | _GEN_312;
    spriteVisibleReg_44 <= reset | _GEN_313;
    spriteVisibleReg_45 <= reset | _GEN_314;
    spriteVisibleReg_46 <= reset | _GEN_315;
    spriteVisibleReg_47 <= reset | _GEN_316;
    spriteVisibleReg_48 <= reset | _GEN_317;
    spriteVisibleReg_49 <= reset | _GEN_318;
    spriteVisibleReg_50 <= reset | _GEN_319;
    spriteVisibleReg_51 <= reset | _GEN_320;
    spriteVisibleReg_55 <= reset | _GEN_324;
    spriteVisibleReg_56 <= reset | _GEN_325;
    spriteVisibleReg_57 <= reset | _GEN_326;
    spriteVisibleReg_61 <= reset | _GEN_330;
    spriteVisibleReg_62 <= reset | _GEN_331;
    spriteVisibleReg_63 <= reset | _GEN_332;
    spriteVisibleReg_64 <= reset | _GEN_333;
    spriteVisibleReg_65 <= reset | _GEN_334;
    spriteVisibleReg_66 <= reset | _GEN_335;
    spriteVisibleReg_70 <= reset | _GEN_339;
    spriteVisibleReg_71 <= reset | _GEN_340;
    spriteVisibleReg_72 <= reset | _GEN_341;
    if (reset) begin
      spriteFlipVerticalReg_122 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_122 <= io_spriteFlipVertical_122;
    end
    if (reset) begin
      spriteFlipVerticalReg_123 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_123 <= io_spriteFlipVertical_123;
    end
    if (reset) begin
      spriteFlipVerticalReg_124 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_124 <= io_spriteFlipVertical_124;
    end
    if (reset) begin
      spriteFlipVerticalReg_125 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_125 <= io_spriteFlipVertical_125;
    end
    if (reset) begin
      spriteFlipVerticalReg_126 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_126 <= io_spriteFlipVertical_126;
    end
    if (reset) begin
      spriteFlipVerticalReg_127 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_127 <= io_spriteFlipVertical_127;
    end
    if (reset) begin
      viewBoxXReg_0 <= 10'h0;
    end else if (io_newFrame) begin
      viewBoxXReg_0 <= io_viewBoxX_0;
    end
    if (reset) begin
      missingFrameErrorReg <= 1'h0;
    end else begin
      missingFrameErrorReg <= _GEN_1172;
    end
    if (reset) begin
      backBufferWriteErrorReg <= 1'h0;
    end else if (_T_415) begin
      backBufferWriteErrorReg <= _GEN_1180;
    end
    if (reset) begin
      viewBoxOutOfRangeErrorReg <= 1'h0;
    end else begin
      viewBoxOutOfRangeErrorReg <= _GEN_1169;
    end
    if (reset) begin
      newFrameStikyReg <= 1'h0;
    end else if (_T_47) begin
      newFrameStikyReg <= 1'h0;
    end else begin
      newFrameStikyReg <= _GEN_1170;
    end
    _T_47 <= io_frameUpdateDone;
    backTileMemoryDataRead_0_0 <= backTileMemories_0_0_io_dataRead;
    backTileMemoryDataRead_0_1 <= backTileMemories_0_1_io_dataRead;
    backTileMemoryDataRead_0_2 <= backTileMemories_0_2_io_dataRead;
    backTileMemoryDataRead_0_3 <= backTileMemories_0_3_io_dataRead;
    backTileMemoryDataRead_0_4 <= backTileMemories_0_4_io_dataRead;
    backTileMemoryDataRead_0_5 <= backTileMemories_0_5_io_dataRead;
    backTileMemoryDataRead_0_6 <= backTileMemories_0_6_io_dataRead;
    backTileMemoryDataRead_0_7 <= backTileMemories_0_7_io_dataRead;
    backTileMemoryDataRead_0_8 <= backTileMemories_0_8_io_dataRead;
    backTileMemoryDataRead_0_9 <= backTileMemories_0_9_io_dataRead;
    backTileMemoryDataRead_0_10 <= backTileMemories_0_10_io_dataRead;
    backTileMemoryDataRead_0_11 <= backTileMemories_0_11_io_dataRead;
    backTileMemoryDataRead_0_12 <= backTileMemories_0_12_io_dataRead;
    backTileMemoryDataRead_0_13 <= backTileMemories_0_13_io_dataRead;
    backTileMemoryDataRead_0_14 <= backTileMemories_0_14_io_dataRead;
    backTileMemoryDataRead_0_15 <= backTileMemories_0_15_io_dataRead;
    backTileMemoryDataRead_0_16 <= backTileMemories_0_16_io_dataRead;
    backTileMemoryDataRead_0_17 <= backTileMemories_0_17_io_dataRead;
    backTileMemoryDataRead_0_18 <= backTileMemories_0_18_io_dataRead;
    backTileMemoryDataRead_0_19 <= backTileMemories_0_19_io_dataRead;
    backTileMemoryDataRead_0_20 <= backTileMemories_0_20_io_dataRead;
    backTileMemoryDataRead_0_21 <= backTileMemories_0_21_io_dataRead;
    backTileMemoryDataRead_0_22 <= backTileMemories_0_22_io_dataRead;
    backTileMemoryDataRead_0_23 <= backTileMemories_0_23_io_dataRead;
    backTileMemoryDataRead_0_24 <= backTileMemories_0_24_io_dataRead;
    backTileMemoryDataRead_0_25 <= backTileMemories_0_25_io_dataRead;
    backTileMemoryDataRead_0_26 <= backTileMemories_0_26_io_dataRead;
    backTileMemoryDataRead_0_27 <= backTileMemories_0_27_io_dataRead;
    backTileMemoryDataRead_0_28 <= backTileMemories_0_28_io_dataRead;
    backTileMemoryDataRead_0_29 <= backTileMemories_0_29_io_dataRead;
    backTileMemoryDataRead_0_30 <= backTileMemories_0_30_io_dataRead;
    backTileMemoryDataRead_0_31 <= backTileMemories_0_31_io_dataRead;
    backTileMemoryDataRead_1_0 <= backTileMemories_1_0_io_dataRead;
    backTileMemoryDataRead_1_1 <= backTileMemories_1_1_io_dataRead;
    backTileMemoryDataRead_1_2 <= backTileMemories_1_2_io_dataRead;
    backTileMemoryDataRead_1_3 <= backTileMemories_1_3_io_dataRead;
    backTileMemoryDataRead_1_4 <= backTileMemories_1_4_io_dataRead;
    backTileMemoryDataRead_1_5 <= backTileMemories_1_5_io_dataRead;
    backTileMemoryDataRead_1_6 <= backTileMemories_1_6_io_dataRead;
    backTileMemoryDataRead_1_7 <= backTileMemories_1_7_io_dataRead;
    backTileMemoryDataRead_1_8 <= backTileMemories_1_8_io_dataRead;
    backTileMemoryDataRead_1_9 <= backTileMemories_1_9_io_dataRead;
    backTileMemoryDataRead_1_10 <= backTileMemories_1_10_io_dataRead;
    backTileMemoryDataRead_1_11 <= backTileMemories_1_11_io_dataRead;
    backTileMemoryDataRead_1_12 <= backTileMemories_1_12_io_dataRead;
    backTileMemoryDataRead_1_13 <= backTileMemories_1_13_io_dataRead;
    backTileMemoryDataRead_1_14 <= backTileMemories_1_14_io_dataRead;
    backTileMemoryDataRead_1_15 <= backTileMemories_1_15_io_dataRead;
    backTileMemoryDataRead_1_16 <= backTileMemories_1_16_io_dataRead;
    backTileMemoryDataRead_1_17 <= backTileMemories_1_17_io_dataRead;
    backTileMemoryDataRead_1_18 <= backTileMemories_1_18_io_dataRead;
    backTileMemoryDataRead_1_19 <= backTileMemories_1_19_io_dataRead;
    backTileMemoryDataRead_1_20 <= backTileMemories_1_20_io_dataRead;
    backTileMemoryDataRead_1_21 <= backTileMemories_1_21_io_dataRead;
    backTileMemoryDataRead_1_22 <= backTileMemories_1_22_io_dataRead;
    backTileMemoryDataRead_1_23 <= backTileMemories_1_23_io_dataRead;
    backTileMemoryDataRead_1_24 <= backTileMemories_1_24_io_dataRead;
    backTileMemoryDataRead_1_25 <= backTileMemories_1_25_io_dataRead;
    backTileMemoryDataRead_1_26 <= backTileMemories_1_26_io_dataRead;
    backTileMemoryDataRead_1_27 <= backTileMemories_1_27_io_dataRead;
    backTileMemoryDataRead_1_28 <= backTileMemories_1_28_io_dataRead;
    backTileMemoryDataRead_1_29 <= backTileMemories_1_29_io_dataRead;
    backTileMemoryDataRead_1_30 <= backTileMemories_1_30_io_dataRead;
    backTileMemoryDataRead_1_31 <= backTileMemories_1_31_io_dataRead;
    if (reset) begin
      backMemoryCopyCounter <= 12'h0;
    end else if (preDisplayArea) begin
      if (_T_369) begin
        backMemoryCopyCounter <= _T_371;
      end
    end else begin
      backMemoryCopyCounter <= 12'h0;
    end
    copyEnabledReg <= preDisplayArea & _T_369;
    _T_377 <= backMemoryRestoreCounter[10:0];
    _T_379 <= io_backBufferWriteAddress;
    _T_382 <= backMemoryRestoreCounter < 12'h800;
    _T_383 <= io_backBufferWriteEnable;
    _T_386 <= io_backBufferWriteData;
    _T_389 <= backMemoryCopyCounter[10:0];
    _T_397 <= backMemoryRestoreCounter[10:0];
    _T_399 <= io_backBufferWriteAddress;
    _T_402 <= backMemoryRestoreCounter < 12'h800;
    _T_403 <= io_backBufferWriteEnable;
    _T_406 <= io_backBufferWriteData;
    _T_409 <= backMemoryCopyCounter[10:0];
    _T_416 <= backBufferMemories_0_io_dataRead;
    _T_419 <= backBufferMemories_1_io_dataRead;
    if (fullBackgroundColor_0[6]) begin
      if (fullBackgroundColor_1[6]) begin
        pixelColorBack <= 6'h0;
      end else begin
        pixelColorBack <= fullBackgroundColor_1[5:0];
      end
    end else begin
      pixelColorBack <= fullBackgroundColor_0[5:0];
    end
    inSpriteX_0 <= $signed(_T_438) - $signed(spriteXPositionReg_0);
    _T_444 <= $signed(_T_442) - $signed(_GEN_1376);
    inSpriteX_1 <= $signed(_T_438) - $signed(spriteXPositionReg_1);
    _T_563 <= $signed(_T_442) - $signed(_GEN_1385);
    inSpriteX_2 <= $signed(_T_438) - $signed(spriteXPositionReg_2);
    _T_682 <= $signed(_T_442) - $signed(_GEN_1394);
    inSpriteX_3 <= $signed(_T_438) - $signed(spriteXPositionReg_3);
    _T_801 <= $signed(_T_442) - $signed(_GEN_1403);
    inSpriteX_4 <= $signed(_T_438) - $signed(spriteXPositionReg_4);
    _T_920 <= $signed(_T_442) - $signed(_GEN_1412);
    inSpriteX_5 <= $signed(_T_438) - $signed(spriteXPositionReg_5);
    _T_1039 <= $signed(_T_442) - $signed(_GEN_1421);
    inSpriteX_6 <= $signed(_T_438) - $signed(spriteXPositionReg_6);
    _T_1158 <= $signed(_T_442) - $signed(_GEN_1430);
    inSpriteX_7 <= $signed(_T_438) - $signed(spriteXPositionReg_7);
    _T_1277 <= $signed(_T_442) - $signed(_GEN_1439);
    inSpriteX_8 <= $signed(_T_438) - $signed(spriteXPositionReg_8);
    _T_1396 <= $signed(_T_442) - $signed(_GEN_1448);
    inSpriteX_9 <= $signed(_T_438) - $signed(spriteXPositionReg_9);
    _T_1515 <= $signed(_T_442) - $signed(_GEN_1457);
    inSpriteX_10 <= $signed(_T_438) - $signed(spriteXPositionReg_10);
    _T_1634 <= $signed(_T_442) - $signed(_GEN_1466);
    inSpriteX_11 <= $signed(_T_438) - $signed(spriteXPositionReg_11);
    _T_1753 <= $signed(_T_442) - $signed(_GEN_1475);
    inSpriteX_12 <= $signed(_T_438) - $signed(spriteXPositionReg_12);
    _T_1872 <= $signed(_T_442) - $signed(_GEN_1484);
    inSpriteX_13 <= $signed(_T_438) - $signed(spriteXPositionReg_13);
    _T_1991 <= $signed(_T_442) - $signed(_GEN_1493);
    inSpriteX_14 <= $signed(_T_438) - $signed(spriteXPositionReg_14);
    _T_2110 <= $signed(_T_442) - $signed(_GEN_1502);
    inSpriteX_15 <= $signed(_T_438) - $signed(spriteXPositionReg_15);
    _T_2229 <= $signed(_T_442) - $signed(_GEN_1511);
    inSpriteX_16 <= $signed(_T_438) - $signed(spriteXPositionReg_16);
    _T_2348 <= $signed(_T_442) - $signed(_GEN_1520);
    inSpriteX_17 <= $signed(_T_438) - $signed(spriteXPositionReg_17);
    _T_2467 <= $signed(_T_442) - $signed(_GEN_1529);
    inSpriteX_18 <= $signed(_T_438) - $signed(spriteXPositionReg_18);
    _T_2586 <= $signed(_T_442) - $signed(_GEN_1538);
    inSpriteX_19 <= $signed(_T_438) - $signed(spriteXPositionReg_19);
    _T_2705 <= $signed(_T_442) - $signed(_GEN_1547);
    inSpriteX_20 <= $signed(_T_438) - $signed(spriteXPositionReg_20);
    _T_2824 <= $signed(_T_442) - $signed(_GEN_1556);
    inSpriteX_21 <= $signed(_T_438) - $signed(spriteXPositionReg_21);
    _T_2943 <= $signed(_T_442) - $signed(_GEN_1565);
    inSpriteX_22 <= $signed(_T_438) - $signed(spriteXPositionReg_22);
    _T_3062 <= $signed(_T_442) - $signed(_GEN_1574);
    inSpriteX_23 <= $signed(_T_438) - $signed(spriteXPositionReg_23);
    _T_3181 <= $signed(_T_442) - $signed(_GEN_1583);
    inSpriteX_24 <= $signed(_T_438) - $signed(spriteXPositionReg_24);
    _T_3300 <= $signed(_T_442) - $signed(_GEN_1592);
    inSpriteX_25 <= $signed(_T_438) - $signed(spriteXPositionReg_25);
    _T_3419 <= $signed(_T_442) - $signed(_GEN_1601);
    inSpriteX_26 <= $signed(_T_438) - $signed(spriteXPositionReg_26);
    _T_3538 <= $signed(_T_442) - $signed(_GEN_1610);
    inSpriteX_27 <= $signed(_T_438) - $signed(spriteXPositionReg_27);
    _T_3657 <= $signed(_T_442) - $signed(_GEN_1619);
    inSpriteX_28 <= $signed(_T_438) - $signed(spriteXPositionReg_28);
    _T_3776 <= $signed(_T_442) - $signed(_GEN_1628);
    inSpriteX_29 <= $signed(_T_438) - $signed(spriteXPositionReg_29);
    _T_3895 <= $signed(_T_442) - $signed(_GEN_1637);
    inSpriteX_30 <= $signed(_T_438) - $signed(spriteXPositionReg_30);
    _T_4014 <= $signed(_T_442) - $signed(_GEN_1646);
    inSpriteX_31 <= $signed(_T_438) - $signed(spriteXPositionReg_31);
    _T_4133 <= $signed(_T_442) - $signed(_GEN_1655);
    inSpriteX_32 <= $signed(_T_438) - $signed(spriteXPositionReg_32);
    _T_4252 <= $signed(_T_442) - $signed(_GEN_1664);
    inSpriteX_33 <= $signed(_T_438) - $signed(spriteXPositionReg_33);
    _T_4371 <= $signed(_T_442) - $signed(_GEN_1673);
    inSpriteX_34 <= $signed(_T_438) - $signed(spriteXPositionReg_34);
    _T_4490 <= $signed(_T_442) - $signed(_GEN_1682);
    inSpriteX_35 <= $signed(_T_438) - $signed(spriteXPositionReg_35);
    _T_4609 <= $signed(_T_442) - $signed(_GEN_1691);
    inSpriteX_36 <= $signed(_T_438) - $signed(spriteXPositionReg_36);
    _T_4728 <= $signed(_T_442) - $signed(_GEN_1700);
    inSpriteX_37 <= $signed(_T_438) - $signed(spriteXPositionReg_37);
    _T_4847 <= $signed(_T_442) - $signed(_GEN_1709);
    inSpriteX_38 <= $signed(_T_438) - $signed(spriteXPositionReg_38);
    _T_4966 <= $signed(_T_442) - $signed(_GEN_1718);
    inSpriteX_39 <= $signed(_T_438) - $signed(spriteXPositionReg_39);
    _T_5085 <= $signed(_T_442) - $signed(_GEN_1727);
    inSpriteX_40 <= $signed(_T_438) - $signed(spriteXPositionReg_40);
    _T_5204 <= $signed(_T_442) - $signed(_GEN_1736);
    inSpriteX_41 <= $signed(_T_438) - $signed(spriteXPositionReg_41);
    _T_5323 <= $signed(_T_442) - $signed(_GEN_1745);
    inSpriteX_42 <= $signed(_T_438) - $signed(spriteXPositionReg_42);
    _T_5442 <= $signed(_T_442) - $signed(_GEN_1754);
    inSpriteX_43 <= $signed(_T_438) - $signed(spriteXPositionReg_43);
    _T_5561 <= $signed(_T_442) - $signed(_GEN_1763);
    inSpriteX_44 <= $signed(_T_438) - $signed(spriteXPositionReg_44);
    _T_5680 <= $signed(_T_442) - $signed(_GEN_1772);
    inSpriteX_45 <= $signed(_T_438) - $signed(spriteXPositionReg_45);
    _T_5799 <= $signed(_T_442) - $signed(_GEN_1781);
    inSpriteX_46 <= $signed(_T_438) - $signed(spriteXPositionReg_46);
    _T_5918 <= $signed(_T_442) - $signed(_GEN_1790);
    inSpriteX_47 <= $signed(_T_438) - $signed(spriteXPositionReg_47);
    _T_6037 <= $signed(_T_442) - $signed(_GEN_1799);
    inSpriteX_48 <= $signed(_T_438) - $signed(spriteXPositionReg_48);
    _T_6156 <= $signed(_T_442) - $signed(_GEN_1808);
    inSpriteX_49 <= $signed(_T_438) - $signed(spriteXPositionReg_49);
    _T_6275 <= $signed(_T_442) - $signed(_GEN_1817);
    inSpriteX_50 <= $signed(_T_438) - $signed(spriteXPositionReg_50);
    _T_6394 <= $signed(_T_442) - $signed(_GEN_1826);
    inSpriteX_51 <= $signed(_T_438) - $signed(spriteXPositionReg_51);
    _T_6513 <= $signed(_T_442) - $signed(_GEN_1835);
    inSpriteX_52 <= $signed(_T_438) - $signed(spriteXPositionReg_52);
    _T_6632 <= $signed(_T_442) - $signed(_GEN_1844);
    inSpriteX_53 <= $signed(_T_438) - $signed(spriteXPositionReg_53);
    _T_6751 <= $signed(_T_442) - $signed(_GEN_1853);
    inSpriteX_54 <= $signed(_T_438) - $signed(spriteXPositionReg_54);
    _T_6870 <= $signed(_T_442) - $signed(_GEN_1862);
    inSpriteX_55 <= $signed(_T_438) - $signed(spriteXPositionReg_55);
    _T_6989 <= $signed(_T_442) - $signed(_GEN_1871);
    inSpriteX_56 <= $signed(_T_438) - $signed(spriteXPositionReg_56);
    _T_7108 <= $signed(_T_442) - $signed(_GEN_1880);
    inSpriteX_57 <= $signed(_T_438) - $signed(spriteXPositionReg_57);
    _T_7227 <= $signed(_T_442) - $signed(_GEN_1889);
    inSpriteX_58 <= $signed(_T_438) - $signed(spriteXPositionReg_58);
    _T_7346 <= $signed(_T_442) - $signed(_GEN_1898);
    inSpriteX_59 <= $signed(_T_438) - $signed(spriteXPositionReg_59);
    _T_7465 <= $signed(_T_442) - $signed(_GEN_1907);
    inSpriteX_60 <= $signed(_T_438) - $signed(spriteXPositionReg_60);
    _T_7584 <= $signed(_T_442) - $signed(_GEN_1916);
    inSpriteX_61 <= $signed(_T_438) - $signed(spriteXPositionReg_61);
    _T_7703 <= $signed(_T_442) - $signed(_GEN_1925);
    inSpriteX_62 <= $signed(_T_438) - $signed(spriteXPositionReg_62);
    _T_7822 <= $signed(_T_442) - $signed(_GEN_1934);
    inSpriteX_63 <= $signed(_T_438) - $signed(spriteXPositionReg_63);
    _T_7941 <= $signed(_T_442) - $signed(_GEN_1943);
    inSpriteX_64 <= $signed(_T_438) - $signed(spriteXPositionReg_64);
    _T_8060 <= $signed(_T_442) - 11'sh0;
    inSpriteX_65 <= $signed(_T_438) - $signed(spriteXPositionReg_65);
    _T_8179 <= $signed(_T_442) - 11'sh0;
    inSpriteX_66 <= $signed(_T_438) - $signed(spriteXPositionReg_66);
    _T_8298 <= $signed(_T_442) - 11'sh0;
    inSpriteX_67 <= $signed(_T_438) - $signed(spriteXPositionReg_67);
    _T_8417 <= $signed(_T_442) - 11'sh0;
    inSpriteX_68 <= $signed(_T_438) - $signed(spriteXPositionReg_68);
    _T_8536 <= $signed(_T_442) - 11'sh0;
    inSpriteX_69 <= $signed(_T_438) - $signed(spriteXPositionReg_69);
    _T_8655 <= $signed(_T_442) - 11'sh0;
    inSpriteX_70 <= $signed(_T_438) - $signed(spriteXPositionReg_70);
    _T_8774 <= $signed(_T_442) - $signed(_GEN_2000);
    inSpriteX_71 <= $signed(_T_438) - $signed(spriteXPositionReg_71);
    _T_8893 <= $signed(_T_442) - $signed(_GEN_2009);
    inSpriteX_72 <= $signed(_T_438) - $signed(spriteXPositionReg_72);
    _T_9012 <= $signed(_T_442) - $signed(_GEN_2018);
    inSpriteX_73 <= $signed(_T_438) - $signed(spriteXPositionReg_73);
    _T_9131 <= $signed(_T_442) - $signed(_GEN_2027);
    inSpriteX_74 <= $signed(_T_438) - $signed(spriteXPositionReg_74);
    _T_9250 <= $signed(_T_442) - $signed(_GEN_2036);
    inSpriteX_75 <= $signed(_T_438) - $signed(spriteXPositionReg_75);
    _T_9369 <= $signed(_T_442) - $signed(_GEN_2045);
    inSpriteX_76 <= $signed(_T_438) - $signed(spriteXPositionReg_76);
    _T_9488 <= $signed(_T_442) - $signed(_GEN_2054);
    inSpriteX_77 <= $signed(_T_438) - $signed(spriteXPositionReg_77);
    _T_9607 <= $signed(_T_442) - $signed(_GEN_2063);
    inSpriteX_78 <= $signed(_T_438) - $signed(spriteXPositionReg_78);
    _T_9726 <= $signed(_T_442) - $signed(_GEN_2072);
    inSpriteX_79 <= $signed(_T_438) - $signed(spriteXPositionReg_79);
    _T_9845 <= $signed(_T_442) - $signed(_GEN_2081);
    inSpriteX_80 <= $signed(_T_438) - $signed(spriteXPositionReg_80);
    _T_9964 <= $signed(_T_442) - $signed(_GEN_2090);
    inSpriteX_81 <= $signed(_T_438) - $signed(spriteXPositionReg_81);
    _T_10083 <= $signed(_T_442) - $signed(_GEN_2099);
    inSpriteX_82 <= $signed(_T_438) - $signed(spriteXPositionReg_82);
    _T_10202 <= $signed(_T_442) - $signed(_GEN_2108);
    inSpriteX_83 <= $signed(_T_438) - $signed(spriteXPositionReg_83);
    _T_10321 <= $signed(_T_442) - $signed(_GEN_2117);
    inSpriteX_84 <= $signed(_T_438) - $signed(spriteXPositionReg_84);
    _T_10440 <= $signed(_T_442) - $signed(_GEN_2126);
    inSpriteX_85 <= $signed(_T_438) - $signed(spriteXPositionReg_85);
    _T_10559 <= $signed(_T_442) - $signed(_GEN_2135);
    inSpriteX_86 <= $signed(_T_438) - $signed(spriteXPositionReg_86);
    _T_10678 <= $signed(_T_442) - $signed(_GEN_2144);
    inSpriteX_87 <= $signed(_T_438) - $signed(spriteXPositionReg_87);
    _T_10797 <= $signed(_T_442) - $signed(_GEN_2153);
    inSpriteX_88 <= $signed(_T_438) - $signed(spriteXPositionReg_88);
    _T_10916 <= $signed(_T_442) - $signed(_GEN_2162);
    inSpriteX_89 <= $signed(_T_438) - $signed(spriteXPositionReg_89);
    _T_11035 <= $signed(_T_442) - $signed(_GEN_2171);
    inSpriteX_90 <= $signed(_T_438) - $signed(spriteXPositionReg_90);
    _T_11154 <= $signed(_T_442) - $signed(_GEN_2180);
    inSpriteX_91 <= $signed(_T_438) - $signed(spriteXPositionReg_91);
    _T_11273 <= $signed(_T_442) - $signed(_GEN_2189);
    inSpriteX_92 <= $signed(_T_438) - $signed(spriteXPositionReg_92);
    _T_11392 <= $signed(_T_442) - $signed(_GEN_2198);
    inSpriteX_93 <= $signed(_T_438) - $signed(spriteXPositionReg_93);
    _T_11511 <= $signed(_T_442) - $signed(_GEN_2207);
    inSpriteX_94 <= $signed(_T_438) - $signed(spriteXPositionReg_94);
    _T_11630 <= $signed(_T_442) - $signed(_GEN_2216);
    inSpriteX_95 <= $signed(_T_438) - $signed(spriteXPositionReg_95);
    _T_11749 <= $signed(_T_442) - $signed(_GEN_2225);
    inSpriteX_96 <= $signed(_T_438) - $signed(spriteXPositionReg_96);
    _T_11868 <= $signed(_T_442) - $signed(_GEN_2234);
    inSpriteX_97 <= $signed(_T_438) - $signed(spriteXPositionReg_97);
    _T_11987 <= $signed(_T_442) - $signed(_GEN_2243);
    inSpriteX_98 <= $signed(_T_438) - $signed(spriteXPositionReg_98);
    _T_12106 <= $signed(_T_442) - $signed(_GEN_2252);
    inSpriteX_99 <= $signed(_T_438) - $signed(spriteXPositionReg_99);
    _T_12225 <= $signed(_T_442) - $signed(_GEN_2261);
    inSpriteX_100 <= $signed(_T_438) - $signed(spriteXPositionReg_100);
    _T_12344 <= $signed(_T_442) - $signed(_GEN_2270);
    inSpriteX_101 <= $signed(_T_438) - $signed(spriteXPositionReg_101);
    _T_12463 <= $signed(_T_442) - $signed(_GEN_2279);
    inSpriteX_102 <= $signed(_T_438) - $signed(spriteXPositionReg_102);
    _T_12582 <= $signed(_T_442) - $signed(_GEN_2288);
    inSpriteX_103 <= $signed(_T_438) - $signed(spriteXPositionReg_103);
    _T_12701 <= $signed(_T_442) - $signed(_GEN_2297);
    inSpriteX_104 <= $signed(_T_438) - $signed(spriteXPositionReg_104);
    _T_12820 <= $signed(_T_442) - $signed(_GEN_2306);
    inSpriteX_105 <= $signed(_T_438) - $signed(spriteXPositionReg_105);
    _T_12939 <= $signed(_T_442) - $signed(_GEN_2315);
    inSpriteX_106 <= $signed(_T_438) - $signed(spriteXPositionReg_106);
    _T_13058 <= $signed(_T_442) - $signed(_GEN_2324);
    inSpriteX_107 <= $signed(_T_438) - $signed(spriteXPositionReg_107);
    _T_13177 <= $signed(_T_442) - $signed(_GEN_2333);
    inSpriteX_108 <= $signed(_T_438) - $signed(spriteXPositionReg_108);
    _T_13296 <= $signed(_T_442) - $signed(_GEN_2342);
    inSpriteX_109 <= $signed(_T_438) - $signed(spriteXPositionReg_109);
    _T_13415 <= $signed(_T_442) - $signed(_GEN_2351);
    inSpriteX_110 <= $signed(_T_438) - $signed(spriteXPositionReg_110);
    _T_13534 <= $signed(_T_442) - $signed(_GEN_2360);
    inSpriteX_111 <= $signed(_T_438) - $signed(spriteXPositionReg_111);
    _T_13653 <= $signed(_T_442) - $signed(_GEN_2369);
    inSpriteX_112 <= $signed(_T_438) - $signed(spriteXPositionReg_112);
    _T_13772 <= $signed(_T_442) - $signed(_GEN_2378);
    inSpriteX_113 <= $signed(_T_438) - $signed(spriteXPositionReg_113);
    _T_13891 <= $signed(_T_442) - $signed(_GEN_2387);
    inSpriteX_114 <= $signed(_T_438) - $signed(spriteXPositionReg_114);
    _T_14010 <= $signed(_T_442) - $signed(_GEN_2396);
    inSpriteX_115 <= $signed(_T_438) - $signed(spriteXPositionReg_115);
    _T_14129 <= $signed(_T_442) - $signed(_GEN_2405);
    inSpriteX_116 <= $signed(_T_438) - $signed(spriteXPositionReg_116);
    _T_14248 <= $signed(_T_442) - $signed(_GEN_2414);
    inSpriteX_117 <= $signed(_T_438) - $signed(spriteXPositionReg_117);
    _T_14367 <= $signed(_T_442) - $signed(_GEN_2423);
    inSpriteX_118 <= $signed(_T_438) - $signed(spriteXPositionReg_118);
    _T_14486 <= $signed(_T_442) - $signed(_GEN_2432);
    inSpriteX_119 <= $signed(_T_438) - $signed(spriteXPositionReg_119);
    _T_14605 <= $signed(_T_442) - $signed(_GEN_2441);
    inSpriteX_120 <= $signed(_T_438) - $signed(spriteXPositionReg_120);
    _T_14724 <= $signed(_T_442) - $signed(_GEN_2450);
    inSpriteX_121 <= $signed(_T_438) - $signed(spriteXPositionReg_121);
    _T_14843 <= $signed(_T_442) - $signed(_GEN_2459);
    inSpriteX_122 <= $signed(_T_438) - $signed(spriteXPositionReg_122);
    _T_14962 <= $signed(_T_442) - $signed(_GEN_2468);
    inSpriteX_123 <= $signed(_T_438) - $signed(spriteXPositionReg_123);
    _T_15081 <= $signed(_T_442) - $signed(_GEN_2477);
    inSpriteX_124 <= $signed(_T_438) - $signed(spriteXPositionReg_124);
    _T_15200 <= $signed(_T_442) - $signed(_GEN_2486);
    inSpriteX_125 <= $signed(_T_438) - $signed(spriteXPositionReg_125);
    _T_15319 <= $signed(_T_442) - $signed(_GEN_2495);
    inSpriteX_126 <= $signed(_T_438) - $signed(spriteXPositionReg_126);
    _T_15438 <= $signed(_T_442) - $signed(_GEN_2504);
    inSpriteX_127 <= $signed(_T_438) - $signed(spriteXPositionReg_127);
    _T_15557 <= $signed(_T_442) - $signed(_GEN_2513);
    _T_15660_0 <= _T_15660_1;
    _T_15660_1 <= _T_15660_2;
    _T_15660_2 <= _T_17 & _T_18;
    _T_15662_0 <= _T_15662_1;
    _T_15662_1 <= _T_15662_2;
    _T_15662_2 <= _T_17 & _T_18;
    _T_15664_0 <= _T_15664_1;
    _T_15664_1 <= _T_15664_2;
    _T_15664_2 <= _T_17 & _T_18;
  end
endmodule
module Memory_326(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_327(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_328(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_329(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_330(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_331(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_332(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_333(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module SoundEngine(
  input        clock,
  input        reset,
  output       io_output_0,
  input  [3:0] io_input
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire  tone_0_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_0_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_0_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_1_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_1_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_1_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_2_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_2_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_2_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_3_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_3_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_3_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_4_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_4_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_4_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_5_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_5_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_5_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_6_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_6_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_6_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_7_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_7_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_7_io_dataRead; // @[SoundEngine.scala 36:23]
  reg  channel_0; // @[SoundEngine.scala 16:30]
  reg  channel_1; // @[SoundEngine.scala 16:30]
  reg  channel_2; // @[SoundEngine.scala 16:30]
  reg  channel_3; // @[SoundEngine.scala 16:30]
  reg  channel_4; // @[SoundEngine.scala 16:30]
  reg  channel_5; // @[SoundEngine.scala 16:30]
  reg  channel_6; // @[SoundEngine.scala 16:30]
  reg  channel_7; // @[SoundEngine.scala 16:30]
  reg [19:0] cntMilliSecond_0; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_1; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_2; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_3; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_4; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_5; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_6; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_7; // @[SoundEngine.scala 17:34]
  reg [19:0] slowCounter_0; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_1; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_2; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_3; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_4; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_5; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_6; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_7; // @[SoundEngine.scala 18:28]
  reg [31:0] waveCnt_0; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_1; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_2; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_3; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_4; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_5; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_6; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_7; // @[SoundEngine.scala 19:28]
  reg [8:0] toneIndex_0; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_1; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_2; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_3; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_4; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_5; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_6; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_7; // @[SoundEngine.scala 20:28]
  reg  songPlaying_0; // @[SoundEngine.scala 21:28]
  reg  songPlaying_1; // @[SoundEngine.scala 21:28]
  reg  songPlaying_2; // @[SoundEngine.scala 21:28]
  reg  songPlaying_3; // @[SoundEngine.scala 21:28]
  reg  songPlaying_4; // @[SoundEngine.scala 21:28]
  reg  songPlaying_5; // @[SoundEngine.scala 21:28]
  reg  songPlaying_6; // @[SoundEngine.scala 21:28]
  reg  songPlaying_7; // @[SoundEngine.scala 21:28]
  wire  _T_9 = io_input > 4'h0; // @[SoundEngine.scala 27:17]
  wire  _T_10 = io_input <= 4'h8; // @[SoundEngine.scala 27:35]
  wire  _T_11 = _T_9 & _T_10; // @[SoundEngine.scala 27:23]
  wire [3:0] _T_13 = io_input - 4'h1; // @[SoundEngine.scala 28:25]
  wire  _GEN_152 = 3'h0 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_8 = _GEN_152 | songPlaying_0; // @[SoundEngine.scala 28:31]
  wire  _GEN_153 = 3'h1 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_9 = _GEN_153 | songPlaying_1; // @[SoundEngine.scala 28:31]
  wire  _GEN_154 = 3'h2 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_10 = _GEN_154 | songPlaying_2; // @[SoundEngine.scala 28:31]
  wire  _GEN_155 = 3'h3 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_11 = _GEN_155 | songPlaying_3; // @[SoundEngine.scala 28:31]
  wire  _GEN_156 = 3'h4 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_12 = _GEN_156 | songPlaying_4; // @[SoundEngine.scala 28:31]
  wire  _GEN_157 = 3'h5 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_13 = _GEN_157 | songPlaying_5; // @[SoundEngine.scala 28:31]
  wire  _GEN_158 = 3'h6 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_14 = _GEN_158 | songPlaying_6; // @[SoundEngine.scala 28:31]
  wire  _GEN_159 = 3'h7 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_15 = _GEN_159 | songPlaying_7; // @[SoundEngine.scala 28:31]
  reg [19:0] freqReg_0; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_1; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_2; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_3; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_4; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_5; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_6; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_7; // @[SoundEngine.scala 49:24]
  reg [11:0] durReg_0; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_1; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_2; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_3; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_4; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_5; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_6; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_7; // @[SoundEngine.scala 50:24]
  wire  _T_39 = ~songPlaying_0; // @[SoundEngine.scala 56:25]
  wire  _T_40 = slowCounter_0 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_42 = cntMilliSecond_0 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_44 = slowCounter_0 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_45 = freqReg_0 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_47 = waveCnt_0 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_160 = {{12'd0}, freqReg_0}; // @[SoundEngine.scala 81:23]
  wire  _T_48 = waveCnt_0 >= _GEN_160; // @[SoundEngine.scala 81:23]
  wire  _T_49 = ~channel_0; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_161 = {{8'd0}, durReg_0}; // @[SoundEngine.scala 88:28]
  wire  _T_50 = cntMilliSecond_0 >= _GEN_161; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_52 = toneIndex_0 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_53 = durReg_0 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_54 = ~songPlaying_1; // @[SoundEngine.scala 56:25]
  wire  _T_55 = slowCounter_1 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_57 = cntMilliSecond_1 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_59 = slowCounter_1 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_60 = freqReg_1 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_62 = waveCnt_1 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_162 = {{12'd0}, freqReg_1}; // @[SoundEngine.scala 81:23]
  wire  _T_63 = waveCnt_1 >= _GEN_162; // @[SoundEngine.scala 81:23]
  wire  _T_64 = ~channel_1; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_163 = {{8'd0}, durReg_1}; // @[SoundEngine.scala 88:28]
  wire  _T_65 = cntMilliSecond_1 >= _GEN_163; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_67 = toneIndex_1 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_68 = durReg_1 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_69 = ~songPlaying_2; // @[SoundEngine.scala 56:25]
  wire  _T_70 = slowCounter_2 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_72 = cntMilliSecond_2 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_74 = slowCounter_2 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_75 = freqReg_2 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_77 = waveCnt_2 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_164 = {{12'd0}, freqReg_2}; // @[SoundEngine.scala 81:23]
  wire  _T_78 = waveCnt_2 >= _GEN_164; // @[SoundEngine.scala 81:23]
  wire  _T_79 = ~channel_2; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_165 = {{8'd0}, durReg_2}; // @[SoundEngine.scala 88:28]
  wire  _T_80 = cntMilliSecond_2 >= _GEN_165; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_82 = toneIndex_2 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_83 = durReg_2 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_84 = ~songPlaying_3; // @[SoundEngine.scala 56:25]
  wire  _T_85 = slowCounter_3 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_87 = cntMilliSecond_3 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_89 = slowCounter_3 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_90 = freqReg_3 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_92 = waveCnt_3 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_166 = {{12'd0}, freqReg_3}; // @[SoundEngine.scala 81:23]
  wire  _T_93 = waveCnt_3 >= _GEN_166; // @[SoundEngine.scala 81:23]
  wire  _T_94 = ~channel_3; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_167 = {{8'd0}, durReg_3}; // @[SoundEngine.scala 88:28]
  wire  _T_95 = cntMilliSecond_3 >= _GEN_167; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_97 = toneIndex_3 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_98 = durReg_3 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_99 = ~songPlaying_4; // @[SoundEngine.scala 56:25]
  wire  _T_100 = slowCounter_4 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_102 = cntMilliSecond_4 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_104 = slowCounter_4 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_105 = freqReg_4 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_107 = waveCnt_4 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_168 = {{12'd0}, freqReg_4}; // @[SoundEngine.scala 81:23]
  wire  _T_108 = waveCnt_4 >= _GEN_168; // @[SoundEngine.scala 81:23]
  wire  _T_109 = ~channel_4; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_169 = {{8'd0}, durReg_4}; // @[SoundEngine.scala 88:28]
  wire  _T_110 = cntMilliSecond_4 >= _GEN_169; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_112 = toneIndex_4 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_113 = durReg_4 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_114 = ~songPlaying_5; // @[SoundEngine.scala 56:25]
  wire  _T_115 = slowCounter_5 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_117 = cntMilliSecond_5 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_119 = slowCounter_5 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_120 = freqReg_5 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_122 = waveCnt_5 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_170 = {{12'd0}, freqReg_5}; // @[SoundEngine.scala 81:23]
  wire  _T_123 = waveCnt_5 >= _GEN_170; // @[SoundEngine.scala 81:23]
  wire  _T_124 = ~channel_5; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_171 = {{8'd0}, durReg_5}; // @[SoundEngine.scala 88:28]
  wire  _T_125 = cntMilliSecond_5 >= _GEN_171; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_127 = toneIndex_5 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_128 = durReg_5 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_129 = ~songPlaying_6; // @[SoundEngine.scala 56:25]
  wire  _T_130 = slowCounter_6 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_132 = cntMilliSecond_6 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_134 = slowCounter_6 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_135 = freqReg_6 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_137 = waveCnt_6 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_172 = {{12'd0}, freqReg_6}; // @[SoundEngine.scala 81:23]
  wire  _T_138 = waveCnt_6 >= _GEN_172; // @[SoundEngine.scala 81:23]
  wire  _T_139 = ~channel_6; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_173 = {{8'd0}, durReg_6}; // @[SoundEngine.scala 88:28]
  wire  _T_140 = cntMilliSecond_6 >= _GEN_173; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_142 = toneIndex_6 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_143 = durReg_6 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_144 = ~songPlaying_7; // @[SoundEngine.scala 56:25]
  wire  _T_145 = slowCounter_7 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_147 = cntMilliSecond_7 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_149 = slowCounter_7 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_150 = freqReg_7 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_152 = waveCnt_7 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_174 = {{12'd0}, freqReg_7}; // @[SoundEngine.scala 81:23]
  wire  _T_153 = waveCnt_7 >= _GEN_174; // @[SoundEngine.scala 81:23]
  wire  _T_154 = ~channel_7; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_175 = {{8'd0}, durReg_7}; // @[SoundEngine.scala 88:28]
  wire  _T_155 = cntMilliSecond_7 >= _GEN_175; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_157 = toneIndex_7 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_158 = durReg_7 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_159 = channel_0 | channel_1; // @[SoundEngine.scala 98:35]
  wire  _T_160 = _T_159 | channel_2; // @[SoundEngine.scala 98:35]
  wire  _T_161 = _T_160 | channel_3; // @[SoundEngine.scala 98:35]
  wire  _T_162 = _T_161 | channel_4; // @[SoundEngine.scala 98:35]
  wire  _T_163 = _T_162 | channel_5; // @[SoundEngine.scala 98:35]
  wire  _T_164 = _T_163 | channel_6; // @[SoundEngine.scala 98:35]
  Memory_326 tone_0 ( // @[SoundEngine.scala 36:23]
    .clock(tone_0_clock),
    .io_address(tone_0_io_address),
    .io_dataRead(tone_0_io_dataRead)
  );
  Memory_327 tone_1 ( // @[SoundEngine.scala 36:23]
    .clock(tone_1_clock),
    .io_address(tone_1_io_address),
    .io_dataRead(tone_1_io_dataRead)
  );
  Memory_328 tone_2 ( // @[SoundEngine.scala 36:23]
    .clock(tone_2_clock),
    .io_address(tone_2_io_address),
    .io_dataRead(tone_2_io_dataRead)
  );
  Memory_329 tone_3 ( // @[SoundEngine.scala 36:23]
    .clock(tone_3_clock),
    .io_address(tone_3_io_address),
    .io_dataRead(tone_3_io_dataRead)
  );
  Memory_330 tone_4 ( // @[SoundEngine.scala 36:23]
    .clock(tone_4_clock),
    .io_address(tone_4_io_address),
    .io_dataRead(tone_4_io_dataRead)
  );
  Memory_331 tone_5 ( // @[SoundEngine.scala 36:23]
    .clock(tone_5_clock),
    .io_address(tone_5_io_address),
    .io_dataRead(tone_5_io_dataRead)
  );
  Memory_332 tone_6 ( // @[SoundEngine.scala 36:23]
    .clock(tone_6_clock),
    .io_address(tone_6_io_address),
    .io_dataRead(tone_6_io_dataRead)
  );
  Memory_333 tone_7 ( // @[SoundEngine.scala 36:23]
    .clock(tone_7_clock),
    .io_address(tone_7_io_address),
    .io_dataRead(tone_7_io_dataRead)
  );
  assign io_output_0 = _T_164 | channel_7; // @[SoundEngine.scala 98:16]
  assign tone_0_clock = clock;
  assign tone_0_io_address = toneIndex_0; // @[SoundEngine.scala 45:24]
  assign tone_1_clock = clock;
  assign tone_1_io_address = toneIndex_1; // @[SoundEngine.scala 45:24]
  assign tone_2_clock = clock;
  assign tone_2_io_address = toneIndex_2; // @[SoundEngine.scala 45:24]
  assign tone_3_clock = clock;
  assign tone_3_io_address = toneIndex_3; // @[SoundEngine.scala 45:24]
  assign tone_4_clock = clock;
  assign tone_4_io_address = toneIndex_4; // @[SoundEngine.scala 45:24]
  assign tone_5_clock = clock;
  assign tone_5_io_address = toneIndex_5; // @[SoundEngine.scala 45:24]
  assign tone_6_clock = clock;
  assign tone_6_io_address = toneIndex_6; // @[SoundEngine.scala 45:24]
  assign tone_7_clock = clock;
  assign tone_7_io_address = toneIndex_7; // @[SoundEngine.scala 45:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  channel_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  channel_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  channel_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  channel_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  channel_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  channel_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  channel_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  channel_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cntMilliSecond_0 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  cntMilliSecond_1 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  cntMilliSecond_2 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  cntMilliSecond_3 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  cntMilliSecond_4 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  cntMilliSecond_5 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  cntMilliSecond_6 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  cntMilliSecond_7 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  slowCounter_0 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  slowCounter_1 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  slowCounter_2 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  slowCounter_3 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  slowCounter_4 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  slowCounter_5 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  slowCounter_6 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  slowCounter_7 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  waveCnt_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  waveCnt_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  waveCnt_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  waveCnt_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  waveCnt_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  waveCnt_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  waveCnt_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  waveCnt_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  toneIndex_0 = _RAND_32[8:0];
  _RAND_33 = {1{`RANDOM}};
  toneIndex_1 = _RAND_33[8:0];
  _RAND_34 = {1{`RANDOM}};
  toneIndex_2 = _RAND_34[8:0];
  _RAND_35 = {1{`RANDOM}};
  toneIndex_3 = _RAND_35[8:0];
  _RAND_36 = {1{`RANDOM}};
  toneIndex_4 = _RAND_36[8:0];
  _RAND_37 = {1{`RANDOM}};
  toneIndex_5 = _RAND_37[8:0];
  _RAND_38 = {1{`RANDOM}};
  toneIndex_6 = _RAND_38[8:0];
  _RAND_39 = {1{`RANDOM}};
  toneIndex_7 = _RAND_39[8:0];
  _RAND_40 = {1{`RANDOM}};
  songPlaying_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  songPlaying_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  songPlaying_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  songPlaying_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  songPlaying_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  songPlaying_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  songPlaying_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  songPlaying_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  freqReg_0 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  freqReg_1 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  freqReg_2 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  freqReg_3 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  freqReg_4 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  freqReg_5 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  freqReg_6 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  freqReg_7 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  durReg_0 = _RAND_56[11:0];
  _RAND_57 = {1{`RANDOM}};
  durReg_1 = _RAND_57[11:0];
  _RAND_58 = {1{`RANDOM}};
  durReg_2 = _RAND_58[11:0];
  _RAND_59 = {1{`RANDOM}};
  durReg_3 = _RAND_59[11:0];
  _RAND_60 = {1{`RANDOM}};
  durReg_4 = _RAND_60[11:0];
  _RAND_61 = {1{`RANDOM}};
  durReg_5 = _RAND_61[11:0];
  _RAND_62 = {1{`RANDOM}};
  durReg_6 = _RAND_62[11:0];
  _RAND_63 = {1{`RANDOM}};
  durReg_7 = _RAND_63[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      channel_0 <= 1'h0;
    end else if (_T_45) begin
      channel_0 <= 1'h0;
    end else if (_T_48) begin
      channel_0 <= _T_49;
    end else if (_T_39) begin
      channel_0 <= 1'h0;
    end
    if (reset) begin
      channel_1 <= 1'h0;
    end else if (_T_60) begin
      channel_1 <= 1'h0;
    end else if (_T_63) begin
      channel_1 <= _T_64;
    end else if (_T_54) begin
      channel_1 <= 1'h0;
    end
    if (reset) begin
      channel_2 <= 1'h0;
    end else if (_T_75) begin
      channel_2 <= 1'h0;
    end else if (_T_78) begin
      channel_2 <= _T_79;
    end else if (_T_69) begin
      channel_2 <= 1'h0;
    end
    if (reset) begin
      channel_3 <= 1'h0;
    end else if (_T_90) begin
      channel_3 <= 1'h0;
    end else if (_T_93) begin
      channel_3 <= _T_94;
    end else if (_T_84) begin
      channel_3 <= 1'h0;
    end
    if (reset) begin
      channel_4 <= 1'h0;
    end else if (_T_105) begin
      channel_4 <= 1'h0;
    end else if (_T_108) begin
      channel_4 <= _T_109;
    end else if (_T_99) begin
      channel_4 <= 1'h0;
    end
    if (reset) begin
      channel_5 <= 1'h0;
    end else if (_T_120) begin
      channel_5 <= 1'h0;
    end else if (_T_123) begin
      channel_5 <= _T_124;
    end else if (_T_114) begin
      channel_5 <= 1'h0;
    end
    if (reset) begin
      channel_6 <= 1'h0;
    end else if (_T_135) begin
      channel_6 <= 1'h0;
    end else if (_T_138) begin
      channel_6 <= _T_139;
    end else if (_T_129) begin
      channel_6 <= 1'h0;
    end
    if (reset) begin
      channel_7 <= 1'h0;
    end else if (_T_150) begin
      channel_7 <= 1'h0;
    end else if (_T_153) begin
      channel_7 <= _T_154;
    end else if (_T_144) begin
      channel_7 <= 1'h0;
    end
    if (reset) begin
      cntMilliSecond_0 <= 20'h0;
    end else if (_T_50) begin
      cntMilliSecond_0 <= 20'h0;
    end else if (_T_40) begin
      cntMilliSecond_0 <= _T_42;
    end else if (_T_39) begin
      cntMilliSecond_0 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_1 <= 20'h0;
    end else if (_T_65) begin
      cntMilliSecond_1 <= 20'h0;
    end else if (_T_55) begin
      cntMilliSecond_1 <= _T_57;
    end else if (_T_54) begin
      cntMilliSecond_1 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_2 <= 20'h0;
    end else if (_T_80) begin
      cntMilliSecond_2 <= 20'h0;
    end else if (_T_70) begin
      cntMilliSecond_2 <= _T_72;
    end else if (_T_69) begin
      cntMilliSecond_2 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_3 <= 20'h0;
    end else if (_T_95) begin
      cntMilliSecond_3 <= 20'h0;
    end else if (_T_85) begin
      cntMilliSecond_3 <= _T_87;
    end else if (_T_84) begin
      cntMilliSecond_3 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_4 <= 20'h0;
    end else if (_T_110) begin
      cntMilliSecond_4 <= 20'h0;
    end else if (_T_100) begin
      cntMilliSecond_4 <= _T_102;
    end else if (_T_99) begin
      cntMilliSecond_4 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_5 <= 20'h0;
    end else if (_T_125) begin
      cntMilliSecond_5 <= 20'h0;
    end else if (_T_115) begin
      cntMilliSecond_5 <= _T_117;
    end else if (_T_114) begin
      cntMilliSecond_5 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_6 <= 20'h0;
    end else if (_T_140) begin
      cntMilliSecond_6 <= 20'h0;
    end else if (_T_130) begin
      cntMilliSecond_6 <= _T_132;
    end else if (_T_129) begin
      cntMilliSecond_6 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_7 <= 20'h0;
    end else if (_T_155) begin
      cntMilliSecond_7 <= 20'h0;
    end else if (_T_145) begin
      cntMilliSecond_7 <= _T_147;
    end else if (_T_144) begin
      cntMilliSecond_7 <= 20'h0;
    end
    if (reset) begin
      slowCounter_0 <= 20'h0;
    end else if (_T_40) begin
      slowCounter_0 <= 20'h0;
    end else begin
      slowCounter_0 <= _T_44;
    end
    if (reset) begin
      slowCounter_1 <= 20'h0;
    end else if (_T_55) begin
      slowCounter_1 <= 20'h0;
    end else begin
      slowCounter_1 <= _T_59;
    end
    if (reset) begin
      slowCounter_2 <= 20'h0;
    end else if (_T_70) begin
      slowCounter_2 <= 20'h0;
    end else begin
      slowCounter_2 <= _T_74;
    end
    if (reset) begin
      slowCounter_3 <= 20'h0;
    end else if (_T_85) begin
      slowCounter_3 <= 20'h0;
    end else begin
      slowCounter_3 <= _T_89;
    end
    if (reset) begin
      slowCounter_4 <= 20'h0;
    end else if (_T_100) begin
      slowCounter_4 <= 20'h0;
    end else begin
      slowCounter_4 <= _T_104;
    end
    if (reset) begin
      slowCounter_5 <= 20'h0;
    end else if (_T_115) begin
      slowCounter_5 <= 20'h0;
    end else begin
      slowCounter_5 <= _T_119;
    end
    if (reset) begin
      slowCounter_6 <= 20'h0;
    end else if (_T_130) begin
      slowCounter_6 <= 20'h0;
    end else begin
      slowCounter_6 <= _T_134;
    end
    if (reset) begin
      slowCounter_7 <= 20'h0;
    end else if (_T_145) begin
      slowCounter_7 <= 20'h0;
    end else begin
      slowCounter_7 <= _T_149;
    end
    if (reset) begin
      waveCnt_0 <= 32'h0;
    end else if (_T_45) begin
      waveCnt_0 <= 32'h0;
    end else if (_T_48) begin
      waveCnt_0 <= 32'h0;
    end else begin
      waveCnt_0 <= _T_47;
    end
    if (reset) begin
      waveCnt_1 <= 32'h0;
    end else if (_T_60) begin
      waveCnt_1 <= 32'h0;
    end else if (_T_63) begin
      waveCnt_1 <= 32'h0;
    end else begin
      waveCnt_1 <= _T_62;
    end
    if (reset) begin
      waveCnt_2 <= 32'h0;
    end else if (_T_75) begin
      waveCnt_2 <= 32'h0;
    end else if (_T_78) begin
      waveCnt_2 <= 32'h0;
    end else begin
      waveCnt_2 <= _T_77;
    end
    if (reset) begin
      waveCnt_3 <= 32'h0;
    end else if (_T_90) begin
      waveCnt_3 <= 32'h0;
    end else if (_T_93) begin
      waveCnt_3 <= 32'h0;
    end else begin
      waveCnt_3 <= _T_92;
    end
    if (reset) begin
      waveCnt_4 <= 32'h0;
    end else if (_T_105) begin
      waveCnt_4 <= 32'h0;
    end else if (_T_108) begin
      waveCnt_4 <= 32'h0;
    end else begin
      waveCnt_4 <= _T_107;
    end
    if (reset) begin
      waveCnt_5 <= 32'h0;
    end else if (_T_120) begin
      waveCnt_5 <= 32'h0;
    end else if (_T_123) begin
      waveCnt_5 <= 32'h0;
    end else begin
      waveCnt_5 <= _T_122;
    end
    if (reset) begin
      waveCnt_6 <= 32'h0;
    end else if (_T_135) begin
      waveCnt_6 <= 32'h0;
    end else if (_T_138) begin
      waveCnt_6 <= 32'h0;
    end else begin
      waveCnt_6 <= _T_137;
    end
    if (reset) begin
      waveCnt_7 <= 32'h0;
    end else if (_T_150) begin
      waveCnt_7 <= 32'h0;
    end else if (_T_153) begin
      waveCnt_7 <= 32'h0;
    end else begin
      waveCnt_7 <= _T_152;
    end
    if (reset) begin
      toneIndex_0 <= 9'h0;
    end else if (_T_50) begin
      toneIndex_0 <= _T_52;
    end else if (_T_39) begin
      toneIndex_0 <= 9'h0;
    end
    if (reset) begin
      toneIndex_1 <= 9'h0;
    end else if (_T_65) begin
      toneIndex_1 <= _T_67;
    end else if (_T_54) begin
      toneIndex_1 <= 9'h0;
    end
    if (reset) begin
      toneIndex_2 <= 9'h0;
    end else if (_T_80) begin
      toneIndex_2 <= _T_82;
    end else if (_T_69) begin
      toneIndex_2 <= 9'h0;
    end
    if (reset) begin
      toneIndex_3 <= 9'h0;
    end else if (_T_95) begin
      toneIndex_3 <= _T_97;
    end else if (_T_84) begin
      toneIndex_3 <= 9'h0;
    end
    if (reset) begin
      toneIndex_4 <= 9'h0;
    end else if (_T_110) begin
      toneIndex_4 <= _T_112;
    end else if (_T_99) begin
      toneIndex_4 <= 9'h0;
    end
    if (reset) begin
      toneIndex_5 <= 9'h0;
    end else if (_T_125) begin
      toneIndex_5 <= _T_127;
    end else if (_T_114) begin
      toneIndex_5 <= 9'h0;
    end
    if (reset) begin
      toneIndex_6 <= 9'h0;
    end else if (_T_140) begin
      toneIndex_6 <= _T_142;
    end else if (_T_129) begin
      toneIndex_6 <= 9'h0;
    end
    if (reset) begin
      toneIndex_7 <= 9'h0;
    end else if (_T_155) begin
      toneIndex_7 <= _T_157;
    end else if (_T_144) begin
      toneIndex_7 <= 9'h0;
    end
    if (reset) begin
      songPlaying_0 <= 1'h0;
    end else if (_T_53) begin
      songPlaying_0 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_0 <= _GEN_8;
    end
    if (reset) begin
      songPlaying_1 <= 1'h0;
    end else if (_T_68) begin
      songPlaying_1 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_1 <= _GEN_9;
    end
    if (reset) begin
      songPlaying_2 <= 1'h0;
    end else if (_T_83) begin
      songPlaying_2 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_2 <= _GEN_10;
    end
    if (reset) begin
      songPlaying_3 <= 1'h0;
    end else if (_T_98) begin
      songPlaying_3 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_3 <= _GEN_11;
    end
    if (reset) begin
      songPlaying_4 <= 1'h0;
    end else if (_T_113) begin
      songPlaying_4 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_4 <= _GEN_12;
    end
    if (reset) begin
      songPlaying_5 <= 1'h0;
    end else if (_T_128) begin
      songPlaying_5 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_5 <= _GEN_13;
    end
    if (reset) begin
      songPlaying_6 <= 1'h0;
    end else if (_T_143) begin
      songPlaying_6 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_6 <= _GEN_14;
    end
    if (reset) begin
      songPlaying_7 <= 1'h0;
    end else if (_T_158) begin
      songPlaying_7 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_7 <= _GEN_15;
    end
    freqReg_0 <= tone_0_io_dataRead[31:12];
    freqReg_1 <= tone_1_io_dataRead[31:12];
    freqReg_2 <= tone_2_io_dataRead[31:12];
    freqReg_3 <= tone_3_io_dataRead[31:12];
    freqReg_4 <= tone_4_io_dataRead[31:12];
    freqReg_5 <= tone_5_io_dataRead[31:12];
    freqReg_6 <= tone_6_io_dataRead[31:12];
    freqReg_7 <= tone_7_io_dataRead[31:12];
    durReg_0 <= tone_0_io_dataRead[11:0];
    durReg_1 <= tone_1_io_dataRead[11:0];
    durReg_2 <= tone_2_io_dataRead[11:0];
    durReg_3 <= tone_3_io_dataRead[11:0];
    durReg_4 <= tone_4_io_dataRead[11:0];
    durReg_5 <= tone_5_io_dataRead[11:0];
    durReg_6 <= tone_6_io_dataRead[11:0];
    durReg_7 <= tone_7_io_dataRead[11:0];
  end
endmodule
module BoxDetection(
  input         clock,
  input  [10:0] io_boxXPosition_0,
  input  [10:0] io_boxXPosition_2,
  input  [10:0] io_boxXPosition_3,
  input  [10:0] io_boxXPosition_4,
  input  [10:0] io_boxXPosition_5,
  input  [10:0] io_boxXPosition_6,
  input  [10:0] io_boxXPosition_7,
  input  [10:0] io_boxXPosition_8,
  input  [10:0] io_boxXPosition_9,
  input  [10:0] io_boxXPosition_10,
  input  [10:0] io_boxXPosition_11,
  input  [10:0] io_boxXPosition_12,
  input  [10:0] io_boxXPosition_13,
  input  [10:0] io_boxXPosition_14,
  input  [10:0] io_boxXPosition_15,
  input  [10:0] io_boxXPosition_16,
  input  [10:0] io_boxXPosition_17,
  input  [9:0]  io_boxYPosition_0,
  input  [9:0]  io_boxYPosition_2,
  input  [9:0]  io_boxYPosition_3,
  input  [9:0]  io_boxYPosition_4,
  input  [9:0]  io_boxYPosition_5,
  input  [9:0]  io_boxYPosition_6,
  input  [9:0]  io_boxYPosition_7,
  input  [9:0]  io_boxYPosition_8,
  input  [9:0]  io_boxYPosition_9,
  input  [9:0]  io_boxYPosition_10,
  input  [9:0]  io_boxYPosition_11,
  input  [9:0]  io_boxYPosition_12,
  input  [9:0]  io_boxYPosition_13,
  input  [9:0]  io_boxYPosition_14,
  input  [9:0]  io_boxYPosition_15,
  input  [9:0]  io_boxYPosition_16,
  input  [9:0]  io_boxYPosition_17,
  output        io_overlap_0_7,
  output        io_overlap_0_8,
  output        io_overlap_0_9,
  output        io_overlap_0_10,
  output        io_overlap_0_11,
  output        io_overlap_0_12,
  output        io_overlap_0_13,
  output        io_overlap_0_14,
  output        io_overlap_0_15,
  output        io_overlap_0_16,
  output        io_overlap_0_17,
  output        io_overlap_2_7,
  output        io_overlap_2_8,
  output        io_overlap_2_9,
  output        io_overlap_2_10,
  output        io_overlap_2_11,
  output        io_overlap_2_12,
  output        io_overlap_2_13,
  output        io_overlap_2_14,
  output        io_overlap_2_15,
  output        io_overlap_2_16,
  output        io_overlap_2_17,
  output        io_overlap_3_7,
  output        io_overlap_3_8,
  output        io_overlap_3_9,
  output        io_overlap_3_10,
  output        io_overlap_3_11,
  output        io_overlap_3_12,
  output        io_overlap_3_13,
  output        io_overlap_3_14,
  output        io_overlap_3_15,
  output        io_overlap_3_16,
  output        io_overlap_3_17,
  output        io_overlap_4_7,
  output        io_overlap_4_8,
  output        io_overlap_4_9,
  output        io_overlap_4_10,
  output        io_overlap_4_11,
  output        io_overlap_4_12,
  output        io_overlap_4_13,
  output        io_overlap_4_14,
  output        io_overlap_4_15,
  output        io_overlap_4_16,
  output        io_overlap_4_17,
  output        io_overlap_5_7,
  output        io_overlap_5_8,
  output        io_overlap_5_9,
  output        io_overlap_5_10,
  output        io_overlap_5_11,
  output        io_overlap_5_12,
  output        io_overlap_5_13,
  output        io_overlap_5_14,
  output        io_overlap_5_15,
  output        io_overlap_5_16,
  output        io_overlap_5_17,
  output        io_overlap_6_7,
  output        io_overlap_6_8,
  output        io_overlap_6_9,
  output        io_overlap_6_10,
  output        io_overlap_6_11,
  output        io_overlap_6_12,
  output        io_overlap_6_13,
  output        io_overlap_6_14,
  output        io_overlap_6_15,
  output        io_overlap_6_17
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  wire [10:0] _T_2 = $signed(io_boxXPosition_0) + 11'sh20; // @[BoxDetection.scala 18:36]
  wire [9:0] _T_5 = $signed(io_boxYPosition_0) + 10'sh20; // @[BoxDetection.scala 19:36]
  wire [10:0] _T_34 = $signed(io_boxXPosition_2) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_37 = $signed(io_boxYPosition_2) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_47 = $signed(io_boxXPosition_3) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_50 = $signed(io_boxYPosition_3) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_60 = $signed(io_boxXPosition_4) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_63 = $signed(io_boxYPosition_4) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_73 = $signed(io_boxXPosition_5) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_76 = $signed(io_boxYPosition_5) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_86 = $signed(io_boxXPosition_6) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_89 = $signed(io_boxYPosition_6) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_99 = $signed(io_boxXPosition_7) + 11'sh8; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_102 = $signed(io_boxYPosition_7) + 10'sh8; // @[BoxDetection.scala 25:38]
  wire  _T_103 = $signed(io_boxXPosition_0) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_104 = $signed(io_boxXPosition_7) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_105 = _T_103 & _T_104; // @[BoxDetection.scala 27:41]
  wire  _T_106 = $signed(io_boxYPosition_0) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_107 = _T_105 & _T_106; // @[BoxDetection.scala 27:60]
  wire  _T_108 = $signed(io_boxYPosition_7) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_112 = $signed(io_boxXPosition_8) + 11'sh10; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_115 = $signed(io_boxYPosition_8) + 10'sh10; // @[BoxDetection.scala 25:38]
  wire  _T_116 = $signed(io_boxXPosition_0) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_117 = $signed(io_boxXPosition_8) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_118 = _T_116 & _T_117; // @[BoxDetection.scala 27:41]
  wire  _T_119 = $signed(io_boxYPosition_0) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_120 = _T_118 & _T_119; // @[BoxDetection.scala 27:60]
  wire  _T_121 = $signed(io_boxYPosition_8) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_125 = $signed(io_boxXPosition_9) + 11'sh1c; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_128 = $signed(io_boxYPosition_9) + 10'sh1c; // @[BoxDetection.scala 25:38]
  wire  _T_129 = $signed(io_boxXPosition_0) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_130 = $signed(io_boxXPosition_9) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_131 = _T_129 & _T_130; // @[BoxDetection.scala 27:41]
  wire  _T_132 = $signed(io_boxYPosition_0) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_133 = _T_131 & _T_132; // @[BoxDetection.scala 27:60]
  wire  _T_134 = $signed(io_boxYPosition_9) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_138 = $signed(io_boxXPosition_10) + 11'sh1c; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_141 = $signed(io_boxYPosition_10) + 10'sh1c; // @[BoxDetection.scala 25:38]
  wire  _T_142 = $signed(io_boxXPosition_0) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_143 = $signed(io_boxXPosition_10) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_144 = _T_142 & _T_143; // @[BoxDetection.scala 27:41]
  wire  _T_145 = $signed(io_boxYPosition_0) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_146 = _T_144 & _T_145; // @[BoxDetection.scala 27:60]
  wire  _T_147 = $signed(io_boxYPosition_10) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_151 = $signed(io_boxXPosition_11) + 11'sh1c; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_154 = $signed(io_boxYPosition_11) + 10'sh1c; // @[BoxDetection.scala 25:38]
  wire  _T_155 = $signed(io_boxXPosition_0) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_156 = $signed(io_boxXPosition_11) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_157 = _T_155 & _T_156; // @[BoxDetection.scala 27:41]
  wire  _T_158 = $signed(io_boxYPosition_0) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_159 = _T_157 & _T_158; // @[BoxDetection.scala 27:60]
  wire  _T_160 = $signed(io_boxYPosition_11) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_164 = $signed(io_boxXPosition_12) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_167 = $signed(io_boxYPosition_12) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_168 = $signed(io_boxXPosition_0) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_169 = $signed(io_boxXPosition_12) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_170 = _T_168 & _T_169; // @[BoxDetection.scala 27:41]
  wire  _T_171 = $signed(io_boxYPosition_0) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_172 = _T_170 & _T_171; // @[BoxDetection.scala 27:60]
  wire  _T_173 = $signed(io_boxYPosition_12) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_177 = $signed(io_boxXPosition_13) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_180 = $signed(io_boxYPosition_13) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_181 = $signed(io_boxXPosition_0) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_182 = $signed(io_boxXPosition_13) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_183 = _T_181 & _T_182; // @[BoxDetection.scala 27:41]
  wire  _T_184 = $signed(io_boxYPosition_0) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_185 = _T_183 & _T_184; // @[BoxDetection.scala 27:60]
  wire  _T_186 = $signed(io_boxYPosition_13) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_190 = $signed(io_boxXPosition_14) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_193 = $signed(io_boxYPosition_14) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_194 = $signed(io_boxXPosition_0) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_195 = $signed(io_boxXPosition_14) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_196 = _T_194 & _T_195; // @[BoxDetection.scala 27:41]
  wire  _T_197 = $signed(io_boxYPosition_0) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_198 = _T_196 & _T_197; // @[BoxDetection.scala 27:60]
  wire  _T_199 = $signed(io_boxYPosition_14) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_203 = $signed(io_boxXPosition_15) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_206 = $signed(io_boxYPosition_15) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_207 = $signed(io_boxXPosition_0) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_208 = $signed(io_boxXPosition_15) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_209 = _T_207 & _T_208; // @[BoxDetection.scala 27:41]
  wire  _T_210 = $signed(io_boxYPosition_0) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_211 = _T_209 & _T_210; // @[BoxDetection.scala 27:60]
  wire  _T_212 = $signed(io_boxYPosition_15) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_216 = $signed(io_boxXPosition_16) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_219 = $signed(io_boxYPosition_16) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_220 = $signed(io_boxXPosition_0) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_221 = $signed(io_boxXPosition_16) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_222 = _T_220 & _T_221; // @[BoxDetection.scala 27:41]
  wire  _T_223 = $signed(io_boxYPosition_0) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_224 = _T_222 & _T_223; // @[BoxDetection.scala 27:60]
  wire  _T_225 = $signed(io_boxYPosition_16) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_229 = $signed(io_boxXPosition_17) + 11'sh60; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_232 = $signed(io_boxYPosition_17) + 10'sh60; // @[BoxDetection.scala 25:38]
  wire  _T_233 = $signed(io_boxXPosition_0) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_234 = $signed(io_boxXPosition_17) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_235 = _T_233 & _T_234; // @[BoxDetection.scala 27:41]
  wire  _T_236 = $signed(io_boxYPosition_0) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_237 = _T_235 & _T_236; // @[BoxDetection.scala 27:60]
  wire  _T_238 = $signed(io_boxYPosition_17) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire  _T_583 = $signed(io_boxXPosition_2) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_584 = $signed(io_boxXPosition_7) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_585 = _T_583 & _T_584; // @[BoxDetection.scala 27:41]
  wire  _T_586 = $signed(io_boxYPosition_2) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_587 = _T_585 & _T_586; // @[BoxDetection.scala 27:60]
  wire  _T_588 = $signed(io_boxYPosition_7) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_596 = $signed(io_boxXPosition_2) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_597 = $signed(io_boxXPosition_8) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_598 = _T_596 & _T_597; // @[BoxDetection.scala 27:41]
  wire  _T_599 = $signed(io_boxYPosition_2) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_600 = _T_598 & _T_599; // @[BoxDetection.scala 27:60]
  wire  _T_601 = $signed(io_boxYPosition_8) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_609 = $signed(io_boxXPosition_2) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_610 = $signed(io_boxXPosition_9) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_611 = _T_609 & _T_610; // @[BoxDetection.scala 27:41]
  wire  _T_612 = $signed(io_boxYPosition_2) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_613 = _T_611 & _T_612; // @[BoxDetection.scala 27:60]
  wire  _T_614 = $signed(io_boxYPosition_9) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_622 = $signed(io_boxXPosition_2) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_623 = $signed(io_boxXPosition_10) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_624 = _T_622 & _T_623; // @[BoxDetection.scala 27:41]
  wire  _T_625 = $signed(io_boxYPosition_2) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_626 = _T_624 & _T_625; // @[BoxDetection.scala 27:60]
  wire  _T_627 = $signed(io_boxYPosition_10) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_635 = $signed(io_boxXPosition_2) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_636 = $signed(io_boxXPosition_11) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_637 = _T_635 & _T_636; // @[BoxDetection.scala 27:41]
  wire  _T_638 = $signed(io_boxYPosition_2) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_639 = _T_637 & _T_638; // @[BoxDetection.scala 27:60]
  wire  _T_640 = $signed(io_boxYPosition_11) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_648 = $signed(io_boxXPosition_2) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_649 = $signed(io_boxXPosition_12) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_650 = _T_648 & _T_649; // @[BoxDetection.scala 27:41]
  wire  _T_651 = $signed(io_boxYPosition_2) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_652 = _T_650 & _T_651; // @[BoxDetection.scala 27:60]
  wire  _T_653 = $signed(io_boxYPosition_12) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_661 = $signed(io_boxXPosition_2) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_662 = $signed(io_boxXPosition_13) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_663 = _T_661 & _T_662; // @[BoxDetection.scala 27:41]
  wire  _T_664 = $signed(io_boxYPosition_2) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_665 = _T_663 & _T_664; // @[BoxDetection.scala 27:60]
  wire  _T_666 = $signed(io_boxYPosition_13) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_674 = $signed(io_boxXPosition_2) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_675 = $signed(io_boxXPosition_14) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_676 = _T_674 & _T_675; // @[BoxDetection.scala 27:41]
  wire  _T_677 = $signed(io_boxYPosition_2) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_678 = _T_676 & _T_677; // @[BoxDetection.scala 27:60]
  wire  _T_679 = $signed(io_boxYPosition_14) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_687 = $signed(io_boxXPosition_2) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_688 = $signed(io_boxXPosition_15) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_689 = _T_687 & _T_688; // @[BoxDetection.scala 27:41]
  wire  _T_690 = $signed(io_boxYPosition_2) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_691 = _T_689 & _T_690; // @[BoxDetection.scala 27:60]
  wire  _T_692 = $signed(io_boxYPosition_15) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_700 = $signed(io_boxXPosition_2) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_701 = $signed(io_boxXPosition_16) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_702 = _T_700 & _T_701; // @[BoxDetection.scala 27:41]
  wire  _T_703 = $signed(io_boxYPosition_2) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_704 = _T_702 & _T_703; // @[BoxDetection.scala 27:60]
  wire  _T_705 = $signed(io_boxYPosition_16) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_713 = $signed(io_boxXPosition_2) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_714 = $signed(io_boxXPosition_17) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_715 = _T_713 & _T_714; // @[BoxDetection.scala 27:41]
  wire  _T_716 = $signed(io_boxYPosition_2) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_717 = _T_715 & _T_716; // @[BoxDetection.scala 27:60]
  wire  _T_718 = $signed(io_boxYPosition_17) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_823 = $signed(io_boxXPosition_3) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_824 = $signed(io_boxXPosition_7) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_825 = _T_823 & _T_824; // @[BoxDetection.scala 27:41]
  wire  _T_826 = $signed(io_boxYPosition_3) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_827 = _T_825 & _T_826; // @[BoxDetection.scala 27:60]
  wire  _T_828 = $signed(io_boxYPosition_7) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_836 = $signed(io_boxXPosition_3) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_837 = $signed(io_boxXPosition_8) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_838 = _T_836 & _T_837; // @[BoxDetection.scala 27:41]
  wire  _T_839 = $signed(io_boxYPosition_3) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_840 = _T_838 & _T_839; // @[BoxDetection.scala 27:60]
  wire  _T_841 = $signed(io_boxYPosition_8) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_849 = $signed(io_boxXPosition_3) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_850 = $signed(io_boxXPosition_9) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_851 = _T_849 & _T_850; // @[BoxDetection.scala 27:41]
  wire  _T_852 = $signed(io_boxYPosition_3) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_853 = _T_851 & _T_852; // @[BoxDetection.scala 27:60]
  wire  _T_854 = $signed(io_boxYPosition_9) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_862 = $signed(io_boxXPosition_3) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_863 = $signed(io_boxXPosition_10) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_864 = _T_862 & _T_863; // @[BoxDetection.scala 27:41]
  wire  _T_865 = $signed(io_boxYPosition_3) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_866 = _T_864 & _T_865; // @[BoxDetection.scala 27:60]
  wire  _T_867 = $signed(io_boxYPosition_10) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_875 = $signed(io_boxXPosition_3) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_876 = $signed(io_boxXPosition_11) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_877 = _T_875 & _T_876; // @[BoxDetection.scala 27:41]
  wire  _T_878 = $signed(io_boxYPosition_3) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_879 = _T_877 & _T_878; // @[BoxDetection.scala 27:60]
  wire  _T_880 = $signed(io_boxYPosition_11) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_888 = $signed(io_boxXPosition_3) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_889 = $signed(io_boxXPosition_12) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_890 = _T_888 & _T_889; // @[BoxDetection.scala 27:41]
  wire  _T_891 = $signed(io_boxYPosition_3) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_892 = _T_890 & _T_891; // @[BoxDetection.scala 27:60]
  wire  _T_893 = $signed(io_boxYPosition_12) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_901 = $signed(io_boxXPosition_3) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_902 = $signed(io_boxXPosition_13) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_903 = _T_901 & _T_902; // @[BoxDetection.scala 27:41]
  wire  _T_904 = $signed(io_boxYPosition_3) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_905 = _T_903 & _T_904; // @[BoxDetection.scala 27:60]
  wire  _T_906 = $signed(io_boxYPosition_13) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_914 = $signed(io_boxXPosition_3) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_915 = $signed(io_boxXPosition_14) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_916 = _T_914 & _T_915; // @[BoxDetection.scala 27:41]
  wire  _T_917 = $signed(io_boxYPosition_3) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_918 = _T_916 & _T_917; // @[BoxDetection.scala 27:60]
  wire  _T_919 = $signed(io_boxYPosition_14) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_927 = $signed(io_boxXPosition_3) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_928 = $signed(io_boxXPosition_15) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_929 = _T_927 & _T_928; // @[BoxDetection.scala 27:41]
  wire  _T_930 = $signed(io_boxYPosition_3) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_931 = _T_929 & _T_930; // @[BoxDetection.scala 27:60]
  wire  _T_932 = $signed(io_boxYPosition_15) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_940 = $signed(io_boxXPosition_3) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_941 = $signed(io_boxXPosition_16) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_942 = _T_940 & _T_941; // @[BoxDetection.scala 27:41]
  wire  _T_943 = $signed(io_boxYPosition_3) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_944 = _T_942 & _T_943; // @[BoxDetection.scala 27:60]
  wire  _T_945 = $signed(io_boxYPosition_16) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_953 = $signed(io_boxXPosition_3) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_954 = $signed(io_boxXPosition_17) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_955 = _T_953 & _T_954; // @[BoxDetection.scala 27:41]
  wire  _T_956 = $signed(io_boxYPosition_3) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_957 = _T_955 & _T_956; // @[BoxDetection.scala 27:60]
  wire  _T_958 = $signed(io_boxYPosition_17) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_1063 = $signed(io_boxXPosition_4) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_1064 = $signed(io_boxXPosition_7) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1065 = _T_1063 & _T_1064; // @[BoxDetection.scala 27:41]
  wire  _T_1066 = $signed(io_boxYPosition_4) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_1067 = _T_1065 & _T_1066; // @[BoxDetection.scala 27:60]
  wire  _T_1068 = $signed(io_boxYPosition_7) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1076 = $signed(io_boxXPosition_4) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_1077 = $signed(io_boxXPosition_8) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1078 = _T_1076 & _T_1077; // @[BoxDetection.scala 27:41]
  wire  _T_1079 = $signed(io_boxYPosition_4) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_1080 = _T_1078 & _T_1079; // @[BoxDetection.scala 27:60]
  wire  _T_1081 = $signed(io_boxYPosition_8) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1089 = $signed(io_boxXPosition_4) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_1090 = $signed(io_boxXPosition_9) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1091 = _T_1089 & _T_1090; // @[BoxDetection.scala 27:41]
  wire  _T_1092 = $signed(io_boxYPosition_4) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_1093 = _T_1091 & _T_1092; // @[BoxDetection.scala 27:60]
  wire  _T_1094 = $signed(io_boxYPosition_9) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1102 = $signed(io_boxXPosition_4) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_1103 = $signed(io_boxXPosition_10) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1104 = _T_1102 & _T_1103; // @[BoxDetection.scala 27:41]
  wire  _T_1105 = $signed(io_boxYPosition_4) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_1106 = _T_1104 & _T_1105; // @[BoxDetection.scala 27:60]
  wire  _T_1107 = $signed(io_boxYPosition_10) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1115 = $signed(io_boxXPosition_4) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_1116 = $signed(io_boxXPosition_11) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1117 = _T_1115 & _T_1116; // @[BoxDetection.scala 27:41]
  wire  _T_1118 = $signed(io_boxYPosition_4) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_1119 = _T_1117 & _T_1118; // @[BoxDetection.scala 27:60]
  wire  _T_1120 = $signed(io_boxYPosition_11) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1128 = $signed(io_boxXPosition_4) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_1129 = $signed(io_boxXPosition_12) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1130 = _T_1128 & _T_1129; // @[BoxDetection.scala 27:41]
  wire  _T_1131 = $signed(io_boxYPosition_4) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_1132 = _T_1130 & _T_1131; // @[BoxDetection.scala 27:60]
  wire  _T_1133 = $signed(io_boxYPosition_12) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1141 = $signed(io_boxXPosition_4) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_1142 = $signed(io_boxXPosition_13) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1143 = _T_1141 & _T_1142; // @[BoxDetection.scala 27:41]
  wire  _T_1144 = $signed(io_boxYPosition_4) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_1145 = _T_1143 & _T_1144; // @[BoxDetection.scala 27:60]
  wire  _T_1146 = $signed(io_boxYPosition_13) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1154 = $signed(io_boxXPosition_4) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_1155 = $signed(io_boxXPosition_14) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1156 = _T_1154 & _T_1155; // @[BoxDetection.scala 27:41]
  wire  _T_1157 = $signed(io_boxYPosition_4) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_1158 = _T_1156 & _T_1157; // @[BoxDetection.scala 27:60]
  wire  _T_1159 = $signed(io_boxYPosition_14) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1167 = $signed(io_boxXPosition_4) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_1168 = $signed(io_boxXPosition_15) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1169 = _T_1167 & _T_1168; // @[BoxDetection.scala 27:41]
  wire  _T_1170 = $signed(io_boxYPosition_4) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_1171 = _T_1169 & _T_1170; // @[BoxDetection.scala 27:60]
  wire  _T_1172 = $signed(io_boxYPosition_15) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1180 = $signed(io_boxXPosition_4) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_1181 = $signed(io_boxXPosition_16) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1182 = _T_1180 & _T_1181; // @[BoxDetection.scala 27:41]
  wire  _T_1183 = $signed(io_boxYPosition_4) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_1184 = _T_1182 & _T_1183; // @[BoxDetection.scala 27:60]
  wire  _T_1185 = $signed(io_boxYPosition_16) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1193 = $signed(io_boxXPosition_4) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_1194 = $signed(io_boxXPosition_17) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1195 = _T_1193 & _T_1194; // @[BoxDetection.scala 27:41]
  wire  _T_1196 = $signed(io_boxYPosition_4) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_1197 = _T_1195 & _T_1196; // @[BoxDetection.scala 27:60]
  wire  _T_1198 = $signed(io_boxYPosition_17) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1303 = $signed(io_boxXPosition_5) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_1304 = $signed(io_boxXPosition_7) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1305 = _T_1303 & _T_1304; // @[BoxDetection.scala 27:41]
  wire  _T_1306 = $signed(io_boxYPosition_5) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_1307 = _T_1305 & _T_1306; // @[BoxDetection.scala 27:60]
  wire  _T_1308 = $signed(io_boxYPosition_7) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1316 = $signed(io_boxXPosition_5) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_1317 = $signed(io_boxXPosition_8) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1318 = _T_1316 & _T_1317; // @[BoxDetection.scala 27:41]
  wire  _T_1319 = $signed(io_boxYPosition_5) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_1320 = _T_1318 & _T_1319; // @[BoxDetection.scala 27:60]
  wire  _T_1321 = $signed(io_boxYPosition_8) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1329 = $signed(io_boxXPosition_5) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_1330 = $signed(io_boxXPosition_9) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1331 = _T_1329 & _T_1330; // @[BoxDetection.scala 27:41]
  wire  _T_1332 = $signed(io_boxYPosition_5) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_1333 = _T_1331 & _T_1332; // @[BoxDetection.scala 27:60]
  wire  _T_1334 = $signed(io_boxYPosition_9) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1342 = $signed(io_boxXPosition_5) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_1343 = $signed(io_boxXPosition_10) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1344 = _T_1342 & _T_1343; // @[BoxDetection.scala 27:41]
  wire  _T_1345 = $signed(io_boxYPosition_5) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_1346 = _T_1344 & _T_1345; // @[BoxDetection.scala 27:60]
  wire  _T_1347 = $signed(io_boxYPosition_10) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1355 = $signed(io_boxXPosition_5) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_1356 = $signed(io_boxXPosition_11) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1357 = _T_1355 & _T_1356; // @[BoxDetection.scala 27:41]
  wire  _T_1358 = $signed(io_boxYPosition_5) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_1359 = _T_1357 & _T_1358; // @[BoxDetection.scala 27:60]
  wire  _T_1360 = $signed(io_boxYPosition_11) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1368 = $signed(io_boxXPosition_5) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_1369 = $signed(io_boxXPosition_12) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1370 = _T_1368 & _T_1369; // @[BoxDetection.scala 27:41]
  wire  _T_1371 = $signed(io_boxYPosition_5) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_1372 = _T_1370 & _T_1371; // @[BoxDetection.scala 27:60]
  wire  _T_1373 = $signed(io_boxYPosition_12) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1381 = $signed(io_boxXPosition_5) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_1382 = $signed(io_boxXPosition_13) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1383 = _T_1381 & _T_1382; // @[BoxDetection.scala 27:41]
  wire  _T_1384 = $signed(io_boxYPosition_5) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_1385 = _T_1383 & _T_1384; // @[BoxDetection.scala 27:60]
  wire  _T_1386 = $signed(io_boxYPosition_13) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1394 = $signed(io_boxXPosition_5) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_1395 = $signed(io_boxXPosition_14) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1396 = _T_1394 & _T_1395; // @[BoxDetection.scala 27:41]
  wire  _T_1397 = $signed(io_boxYPosition_5) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_1398 = _T_1396 & _T_1397; // @[BoxDetection.scala 27:60]
  wire  _T_1399 = $signed(io_boxYPosition_14) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1407 = $signed(io_boxXPosition_5) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_1408 = $signed(io_boxXPosition_15) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1409 = _T_1407 & _T_1408; // @[BoxDetection.scala 27:41]
  wire  _T_1410 = $signed(io_boxYPosition_5) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_1411 = _T_1409 & _T_1410; // @[BoxDetection.scala 27:60]
  wire  _T_1412 = $signed(io_boxYPosition_15) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1420 = $signed(io_boxXPosition_5) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_1421 = $signed(io_boxXPosition_16) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1422 = _T_1420 & _T_1421; // @[BoxDetection.scala 27:41]
  wire  _T_1423 = $signed(io_boxYPosition_5) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_1424 = _T_1422 & _T_1423; // @[BoxDetection.scala 27:60]
  wire  _T_1425 = $signed(io_boxYPosition_16) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1433 = $signed(io_boxXPosition_5) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_1434 = $signed(io_boxXPosition_17) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1435 = _T_1433 & _T_1434; // @[BoxDetection.scala 27:41]
  wire  _T_1436 = $signed(io_boxYPosition_5) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_1437 = _T_1435 & _T_1436; // @[BoxDetection.scala 27:60]
  wire  _T_1438 = $signed(io_boxYPosition_17) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1543 = $signed(io_boxXPosition_6) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_1544 = $signed(io_boxXPosition_7) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1545 = _T_1543 & _T_1544; // @[BoxDetection.scala 27:41]
  wire  _T_1546 = $signed(io_boxYPosition_6) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_1547 = _T_1545 & _T_1546; // @[BoxDetection.scala 27:60]
  wire  _T_1548 = $signed(io_boxYPosition_7) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1556 = $signed(io_boxXPosition_6) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_1557 = $signed(io_boxXPosition_8) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1558 = _T_1556 & _T_1557; // @[BoxDetection.scala 27:41]
  wire  _T_1559 = $signed(io_boxYPosition_6) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_1560 = _T_1558 & _T_1559; // @[BoxDetection.scala 27:60]
  wire  _T_1561 = $signed(io_boxYPosition_8) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1569 = $signed(io_boxXPosition_6) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_1570 = $signed(io_boxXPosition_9) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1571 = _T_1569 & _T_1570; // @[BoxDetection.scala 27:41]
  wire  _T_1572 = $signed(io_boxYPosition_6) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_1573 = _T_1571 & _T_1572; // @[BoxDetection.scala 27:60]
  wire  _T_1574 = $signed(io_boxYPosition_9) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1582 = $signed(io_boxXPosition_6) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_1583 = $signed(io_boxXPosition_10) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1584 = _T_1582 & _T_1583; // @[BoxDetection.scala 27:41]
  wire  _T_1585 = $signed(io_boxYPosition_6) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_1586 = _T_1584 & _T_1585; // @[BoxDetection.scala 27:60]
  wire  _T_1587 = $signed(io_boxYPosition_10) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1595 = $signed(io_boxXPosition_6) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_1596 = $signed(io_boxXPosition_11) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1597 = _T_1595 & _T_1596; // @[BoxDetection.scala 27:41]
  wire  _T_1598 = $signed(io_boxYPosition_6) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_1599 = _T_1597 & _T_1598; // @[BoxDetection.scala 27:60]
  wire  _T_1600 = $signed(io_boxYPosition_11) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1608 = $signed(io_boxXPosition_6) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_1609 = $signed(io_boxXPosition_12) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1610 = _T_1608 & _T_1609; // @[BoxDetection.scala 27:41]
  wire  _T_1611 = $signed(io_boxYPosition_6) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_1612 = _T_1610 & _T_1611; // @[BoxDetection.scala 27:60]
  wire  _T_1613 = $signed(io_boxYPosition_12) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1621 = $signed(io_boxXPosition_6) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_1622 = $signed(io_boxXPosition_13) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1623 = _T_1621 & _T_1622; // @[BoxDetection.scala 27:41]
  wire  _T_1624 = $signed(io_boxYPosition_6) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_1625 = _T_1623 & _T_1624; // @[BoxDetection.scala 27:60]
  wire  _T_1626 = $signed(io_boxYPosition_13) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1634 = $signed(io_boxXPosition_6) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_1635 = $signed(io_boxXPosition_14) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1636 = _T_1634 & _T_1635; // @[BoxDetection.scala 27:41]
  wire  _T_1637 = $signed(io_boxYPosition_6) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_1638 = _T_1636 & _T_1637; // @[BoxDetection.scala 27:60]
  wire  _T_1639 = $signed(io_boxYPosition_14) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1647 = $signed(io_boxXPosition_6) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_1648 = $signed(io_boxXPosition_15) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1649 = _T_1647 & _T_1648; // @[BoxDetection.scala 27:41]
  wire  _T_1650 = $signed(io_boxYPosition_6) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_1651 = _T_1649 & _T_1650; // @[BoxDetection.scala 27:60]
  wire  _T_1652 = $signed(io_boxYPosition_15) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1673 = $signed(io_boxXPosition_6) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_1674 = $signed(io_boxXPosition_17) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1675 = _T_1673 & _T_1674; // @[BoxDetection.scala 27:41]
  wire  _T_1676 = $signed(io_boxYPosition_6) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_1677 = _T_1675 & _T_1676; // @[BoxDetection.scala 27:60]
  wire  _T_1678 = $signed(io_boxYPosition_17) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  reg  _T_4320_0_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_17; // @[BoxDetection.scala 32:24]
  assign io_overlap_0_7 = _T_4320_0_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_8 = _T_4320_0_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_9 = _T_4320_0_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_10 = _T_4320_0_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_11 = _T_4320_0_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_12 = _T_4320_0_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_13 = _T_4320_0_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_14 = _T_4320_0_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_15 = _T_4320_0_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_16 = _T_4320_0_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_17 = _T_4320_0_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_7 = _T_4320_2_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_8 = _T_4320_2_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_9 = _T_4320_2_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_10 = _T_4320_2_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_11 = _T_4320_2_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_12 = _T_4320_2_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_13 = _T_4320_2_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_14 = _T_4320_2_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_15 = _T_4320_2_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_16 = _T_4320_2_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_17 = _T_4320_2_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_7 = _T_4320_3_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_8 = _T_4320_3_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_9 = _T_4320_3_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_10 = _T_4320_3_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_11 = _T_4320_3_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_12 = _T_4320_3_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_13 = _T_4320_3_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_14 = _T_4320_3_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_15 = _T_4320_3_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_16 = _T_4320_3_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_17 = _T_4320_3_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_7 = _T_4320_4_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_8 = _T_4320_4_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_9 = _T_4320_4_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_10 = _T_4320_4_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_11 = _T_4320_4_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_12 = _T_4320_4_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_13 = _T_4320_4_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_14 = _T_4320_4_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_15 = _T_4320_4_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_16 = _T_4320_4_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_17 = _T_4320_4_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_7 = _T_4320_5_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_8 = _T_4320_5_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_9 = _T_4320_5_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_10 = _T_4320_5_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_11 = _T_4320_5_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_12 = _T_4320_5_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_13 = _T_4320_5_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_14 = _T_4320_5_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_15 = _T_4320_5_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_16 = _T_4320_5_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_17 = _T_4320_5_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_7 = _T_4320_6_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_8 = _T_4320_6_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_9 = _T_4320_6_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_10 = _T_4320_6_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_11 = _T_4320_6_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_12 = _T_4320_6_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_13 = _T_4320_6_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_14 = _T_4320_6_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_15 = _T_4320_6_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_17 = _T_4320_6_17; // @[BoxDetection.scala 32:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4320_0_7 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_4320_0_8 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_4320_0_9 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_4320_0_10 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_4320_0_11 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_4320_0_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_4320_0_13 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_4320_0_14 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_4320_0_15 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_4320_0_16 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_4320_0_17 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_4320_2_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_4320_2_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_4320_2_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_4320_2_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_4320_2_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_4320_2_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_4320_2_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_4320_2_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_4320_2_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_4320_2_16 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4320_2_17 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4320_3_7 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4320_3_8 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4320_3_9 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4320_3_10 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4320_3_11 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4320_3_12 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4320_3_13 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4320_3_14 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4320_3_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4320_3_16 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4320_3_17 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4320_4_7 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4320_4_8 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4320_4_9 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4320_4_10 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4320_4_11 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4320_4_12 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4320_4_13 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4320_4_14 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4320_4_15 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4320_4_16 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4320_4_17 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4320_5_7 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4320_5_8 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4320_5_9 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4320_5_10 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4320_5_11 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4320_5_12 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4320_5_13 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4320_5_14 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4320_5_15 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4320_5_16 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4320_5_17 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4320_6_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4320_6_8 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4320_6_9 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4320_6_10 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4320_6_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4320_6_12 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4320_6_13 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4320_6_14 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4320_6_15 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4320_6_17 = _RAND_64[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_4320_0_7 <= _T_107 & _T_108;
    _T_4320_0_8 <= _T_120 & _T_121;
    _T_4320_0_9 <= _T_133 & _T_134;
    _T_4320_0_10 <= _T_146 & _T_147;
    _T_4320_0_11 <= _T_159 & _T_160;
    _T_4320_0_12 <= _T_172 & _T_173;
    _T_4320_0_13 <= _T_185 & _T_186;
    _T_4320_0_14 <= _T_198 & _T_199;
    _T_4320_0_15 <= _T_211 & _T_212;
    _T_4320_0_16 <= _T_224 & _T_225;
    _T_4320_0_17 <= _T_237 & _T_238;
    _T_4320_2_7 <= _T_587 & _T_588;
    _T_4320_2_8 <= _T_600 & _T_601;
    _T_4320_2_9 <= _T_613 & _T_614;
    _T_4320_2_10 <= _T_626 & _T_627;
    _T_4320_2_11 <= _T_639 & _T_640;
    _T_4320_2_12 <= _T_652 & _T_653;
    _T_4320_2_13 <= _T_665 & _T_666;
    _T_4320_2_14 <= _T_678 & _T_679;
    _T_4320_2_15 <= _T_691 & _T_692;
    _T_4320_2_16 <= _T_704 & _T_705;
    _T_4320_2_17 <= _T_717 & _T_718;
    _T_4320_3_7 <= _T_827 & _T_828;
    _T_4320_3_8 <= _T_840 & _T_841;
    _T_4320_3_9 <= _T_853 & _T_854;
    _T_4320_3_10 <= _T_866 & _T_867;
    _T_4320_3_11 <= _T_879 & _T_880;
    _T_4320_3_12 <= _T_892 & _T_893;
    _T_4320_3_13 <= _T_905 & _T_906;
    _T_4320_3_14 <= _T_918 & _T_919;
    _T_4320_3_15 <= _T_931 & _T_932;
    _T_4320_3_16 <= _T_944 & _T_945;
    _T_4320_3_17 <= _T_957 & _T_958;
    _T_4320_4_7 <= _T_1067 & _T_1068;
    _T_4320_4_8 <= _T_1080 & _T_1081;
    _T_4320_4_9 <= _T_1093 & _T_1094;
    _T_4320_4_10 <= _T_1106 & _T_1107;
    _T_4320_4_11 <= _T_1119 & _T_1120;
    _T_4320_4_12 <= _T_1132 & _T_1133;
    _T_4320_4_13 <= _T_1145 & _T_1146;
    _T_4320_4_14 <= _T_1158 & _T_1159;
    _T_4320_4_15 <= _T_1171 & _T_1172;
    _T_4320_4_16 <= _T_1184 & _T_1185;
    _T_4320_4_17 <= _T_1197 & _T_1198;
    _T_4320_5_7 <= _T_1307 & _T_1308;
    _T_4320_5_8 <= _T_1320 & _T_1321;
    _T_4320_5_9 <= _T_1333 & _T_1334;
    _T_4320_5_10 <= _T_1346 & _T_1347;
    _T_4320_5_11 <= _T_1359 & _T_1360;
    _T_4320_5_12 <= _T_1372 & _T_1373;
    _T_4320_5_13 <= _T_1385 & _T_1386;
    _T_4320_5_14 <= _T_1398 & _T_1399;
    _T_4320_5_15 <= _T_1411 & _T_1412;
    _T_4320_5_16 <= _T_1424 & _T_1425;
    _T_4320_5_17 <= _T_1437 & _T_1438;
    _T_4320_6_7 <= _T_1547 & _T_1548;
    _T_4320_6_8 <= _T_1560 & _T_1561;
    _T_4320_6_9 <= _T_1573 & _T_1574;
    _T_4320_6_10 <= _T_1586 & _T_1587;
    _T_4320_6_11 <= _T_1599 & _T_1600;
    _T_4320_6_12 <= _T_1612 & _T_1613;
    _T_4320_6_13 <= _T_1625 & _T_1626;
    _T_4320_6_14 <= _T_1638 & _T_1639;
    _T_4320_6_15 <= _T_1651 & _T_1652;
    _T_4320_6_17 <= _T_1677 & _T_1678;
  end
endmodule
module Randomizer(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_1(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_2(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h8;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_3(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h8;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_4(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h9;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_5(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h9;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_6(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'ha;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_7(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'ha;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_8(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hb;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_9(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hb;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_10(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hc;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_11(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hc;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_12(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hd;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_13(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hd;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_14(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'he;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_15(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'he;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_16(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hf;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_17(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hf;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_18(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h10;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_19(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h10;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_33(
  input        clock,
  input        reset,
  output [1:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [1:0] place; // @[Randomizer.scala 19:22]
  reg [1:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 2'h2; // @[Randomizer.scala 26:14]
  wire [2:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h1;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 2'h0;
    end else begin
      place <= {{1'd0}, state[0]};
    end
    if (reset) begin
      placeholder <= 2'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[1:0];
    end
  end
endmodule
module Randomizer_34(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7d;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_35(
  input        clock,
  input        reset,
  output [5:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [5:0] place; // @[Randomizer.scala 19:22]
  reg [5:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 6'h11; // @[Randomizer.scala 26:14]
  wire [6:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h9;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 6'h0;
    end else begin
      place <= {{1'd0}, state[4:0]};
    end
    if (reset) begin
      placeholder <= 6'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[5:0];
    end
  end
endmodule
module Randomizer_36(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7e;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_38(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7f;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_40(
  input        clock,
  input        reset,
  output [1:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [1:0] place; // @[Randomizer.scala 19:22]
  reg [1:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 2'h2; // @[Randomizer.scala 26:14]
  wire [2:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h2;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 2'h0;
    end else begin
      place <= {{1'd0}, state[0]};
    end
    if (reset) begin
      placeholder <= 2'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[1:0];
    end
  end
endmodule
module Randomizer_41(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7a;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_43(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7b;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_45(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7c;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module GameLogic(
  input         clock,
  input         reset,
  input         io_btnC,
  input         io_btnU,
  input         io_btnL,
  input         io_btnR,
  input         io_btnD,
  input         io_sw_0,
  input         io_sw_1,
  input         io_sw_2,
  input         io_sw_7,
  output [3:0]  io_songInput,
  output [10:0] io_spriteXPosition_0,
  output [10:0] io_spriteXPosition_1,
  output [10:0] io_spriteXPosition_2,
  output [10:0] io_spriteXPosition_3,
  output [10:0] io_spriteXPosition_4,
  output [10:0] io_spriteXPosition_5,
  output [10:0] io_spriteXPosition_6,
  output [10:0] io_spriteXPosition_7,
  output [10:0] io_spriteXPosition_8,
  output [10:0] io_spriteXPosition_9,
  output [10:0] io_spriteXPosition_10,
  output [10:0] io_spriteXPosition_11,
  output [10:0] io_spriteXPosition_12,
  output [10:0] io_spriteXPosition_13,
  output [10:0] io_spriteXPosition_14,
  output [10:0] io_spriteXPosition_15,
  output [10:0] io_spriteXPosition_16,
  output [10:0] io_spriteXPosition_17,
  output [10:0] io_spriteXPosition_18,
  output [10:0] io_spriteXPosition_19,
  output [10:0] io_spriteXPosition_20,
  output [10:0] io_spriteXPosition_21,
  output [10:0] io_spriteXPosition_22,
  output [10:0] io_spriteXPosition_23,
  output [10:0] io_spriteXPosition_24,
  output [10:0] io_spriteXPosition_25,
  output [10:0] io_spriteXPosition_26,
  output [10:0] io_spriteXPosition_27,
  output [10:0] io_spriteXPosition_28,
  output [10:0] io_spriteXPosition_29,
  output [10:0] io_spriteXPosition_30,
  output [10:0] io_spriteXPosition_31,
  output [10:0] io_spriteXPosition_32,
  output [10:0] io_spriteXPosition_33,
  output [10:0] io_spriteXPosition_41,
  output [10:0] io_spriteXPosition_42,
  output [10:0] io_spriteXPosition_43,
  output [10:0] io_spriteXPosition_44,
  output [10:0] io_spriteXPosition_45,
  output [10:0] io_spriteXPosition_46,
  output [10:0] io_spriteXPosition_47,
  output [10:0] io_spriteXPosition_48,
  output [10:0] io_spriteXPosition_49,
  output [10:0] io_spriteXPosition_50,
  output [10:0] io_spriteXPosition_51,
  output [10:0] io_spriteXPosition_122,
  output [10:0] io_spriteXPosition_123,
  output [10:0] io_spriteXPosition_124,
  output [10:0] io_spriteXPosition_125,
  output [10:0] io_spriteXPosition_126,
  output [10:0] io_spriteXPosition_127,
  output [9:0]  io_spriteYPosition_0,
  output [9:0]  io_spriteYPosition_1,
  output [9:0]  io_spriteYPosition_2,
  output [9:0]  io_spriteYPosition_3,
  output [9:0]  io_spriteYPosition_4,
  output [9:0]  io_spriteYPosition_5,
  output [9:0]  io_spriteYPosition_6,
  output [9:0]  io_spriteYPosition_7,
  output [9:0]  io_spriteYPosition_8,
  output [9:0]  io_spriteYPosition_9,
  output [9:0]  io_spriteYPosition_10,
  output [9:0]  io_spriteYPosition_11,
  output [9:0]  io_spriteYPosition_12,
  output [9:0]  io_spriteYPosition_13,
  output [9:0]  io_spriteYPosition_14,
  output [9:0]  io_spriteYPosition_15,
  output [9:0]  io_spriteYPosition_16,
  output [9:0]  io_spriteYPosition_17,
  output [9:0]  io_spriteYPosition_18,
  output [9:0]  io_spriteYPosition_19,
  output [9:0]  io_spriteYPosition_20,
  output [9:0]  io_spriteYPosition_21,
  output [9:0]  io_spriteYPosition_22,
  output [9:0]  io_spriteYPosition_23,
  output [9:0]  io_spriteYPosition_24,
  output [9:0]  io_spriteYPosition_25,
  output [9:0]  io_spriteYPosition_26,
  output [9:0]  io_spriteYPosition_27,
  output [9:0]  io_spriteYPosition_28,
  output [9:0]  io_spriteYPosition_29,
  output [9:0]  io_spriteYPosition_30,
  output [9:0]  io_spriteYPosition_31,
  output [9:0]  io_spriteYPosition_32,
  output [9:0]  io_spriteYPosition_33,
  output [9:0]  io_spriteYPosition_41,
  output [9:0]  io_spriteYPosition_42,
  output [9:0]  io_spriteYPosition_43,
  output [9:0]  io_spriteYPosition_122,
  output [9:0]  io_spriteYPosition_123,
  output [9:0]  io_spriteYPosition_124,
  output [9:0]  io_spriteYPosition_125,
  output [9:0]  io_spriteYPosition_126,
  output [9:0]  io_spriteYPosition_127,
  output        io_spriteVisible_0,
  output        io_spriteVisible_1,
  output        io_spriteVisible_2,
  output        io_spriteVisible_3,
  output        io_spriteVisible_4,
  output        io_spriteVisible_5,
  output        io_spriteVisible_6,
  output        io_spriteVisible_7,
  output        io_spriteVisible_8,
  output        io_spriteVisible_9,
  output        io_spriteVisible_10,
  output        io_spriteVisible_11,
  output        io_spriteVisible_12,
  output        io_spriteVisible_13,
  output        io_spriteVisible_14,
  output        io_spriteVisible_15,
  output        io_spriteVisible_16,
  output        io_spriteVisible_17,
  output        io_spriteVisible_18,
  output        io_spriteVisible_19,
  output        io_spriteVisible_20,
  output        io_spriteVisible_21,
  output        io_spriteVisible_22,
  output        io_spriteVisible_23,
  output        io_spriteVisible_24,
  output        io_spriteVisible_25,
  output        io_spriteVisible_26,
  output        io_spriteVisible_27,
  output        io_spriteVisible_28,
  output        io_spriteVisible_29,
  output        io_spriteVisible_30,
  output        io_spriteVisible_31,
  output        io_spriteVisible_32,
  output        io_spriteVisible_33,
  output        io_spriteVisible_41,
  output        io_spriteVisible_42,
  output        io_spriteVisible_43,
  output        io_spriteVisible_44,
  output        io_spriteVisible_45,
  output        io_spriteVisible_46,
  output        io_spriteVisible_47,
  output        io_spriteVisible_48,
  output        io_spriteVisible_49,
  output        io_spriteVisible_50,
  output        io_spriteVisible_51,
  output        io_spriteVisible_55,
  output        io_spriteVisible_56,
  output        io_spriteVisible_57,
  output        io_spriteVisible_61,
  output        io_spriteVisible_62,
  output        io_spriteVisible_63,
  output        io_spriteVisible_64,
  output        io_spriteVisible_65,
  output        io_spriteVisible_66,
  output        io_spriteVisible_70,
  output        io_spriteVisible_71,
  output        io_spriteVisible_72,
  output        io_spriteFlipVertical_122,
  output        io_spriteFlipVertical_123,
  output        io_spriteFlipVertical_124,
  output        io_spriteFlipVertical_125,
  output        io_spriteFlipVertical_126,
  output        io_spriteFlipVertical_127,
  output [9:0]  io_viewBoxX_0,
  output [4:0]  io_backBufferWriteData,
  output [10:0] io_backBufferWriteAddress,
  output        io_backBufferWriteEnable,
  input         io_newFrame,
  output        io_frameUpdateDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
`endif // RANDOMIZE_REG_INIT
  wire  boxDetection_clock; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_0; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_2; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_3; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_4; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_5; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_6; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_7; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_8; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_9; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_10; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_11; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_12; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_13; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_14; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_15; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_16; // @[GameLogic.scala 712:28]
  wire [10:0] boxDetection_io_boxXPosition_17; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_0; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_2; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_3; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_4; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_5; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_6; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_7; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_8; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_9; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_10; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_11; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_12; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_13; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_14; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_15; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_16; // @[GameLogic.scala 712:28]
  wire [9:0] boxDetection_io_boxYPosition_17; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_7; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_8; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_9; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_10; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_11; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_12; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_13; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_14; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_15; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_16; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_0_17; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_7; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_8; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_9; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_10; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_11; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_12; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_13; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_14; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_15; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_16; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_2_17; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_7; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_8; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_9; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_10; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_11; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_12; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_13; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_14; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_15; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_16; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_3_17; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_7; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_8; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_9; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_10; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_11; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_12; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_13; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_14; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_15; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_16; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_4_17; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_7; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_8; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_9; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_10; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_11; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_12; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_13; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_14; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_15; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_16; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_5_17; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_7; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_8; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_9; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_10; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_11; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_12; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_13; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_14; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_15; // @[GameLogic.scala 712:28]
  wire  boxDetection_io_overlap_6_17; // @[GameLogic.scala 712:28]
  wire  Randomizer_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_1_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_1_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_1_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_2_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_2_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_2_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_3_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_3_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_3_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_4_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_4_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_4_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_5_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_5_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_5_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_6_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_6_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_6_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_7_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_7_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_7_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_8_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_8_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_8_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_9_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_9_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_9_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_10_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_10_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_10_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_11_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_11_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_11_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_12_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_12_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_12_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_13_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_13_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_13_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_14_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_14_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_14_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_15_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_15_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_15_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_16_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_16_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_16_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_17_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_17_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_17_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_18_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_18_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_18_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_19_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_19_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_19_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_20_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_20_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_20_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_21_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_21_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_21_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_22_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_22_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_22_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_23_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_23_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_23_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_24_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_24_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_24_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_25_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_25_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_25_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_26_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_26_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_26_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_27_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_27_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_27_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_28_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_28_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_28_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_29_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_29_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_29_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_30_clock; // @[GameLogic.scala 201:24]
  wire  Randomizer_30_reset; // @[GameLogic.scala 201:24]
  wire [9:0] Randomizer_30_io_out; // @[GameLogic.scala 201:24]
  wire  Randomizer_31_clock; // @[GameLogic.scala 202:31]
  wire  Randomizer_31_reset; // @[GameLogic.scala 202:31]
  wire [6:0] Randomizer_31_io_out; // @[GameLogic.scala 202:31]
  wire  Randomizer_32_clock; // @[GameLogic.scala 374:24]
  wire  Randomizer_32_reset; // @[GameLogic.scala 374:24]
  wire [9:0] Randomizer_32_io_out; // @[GameLogic.scala 374:24]
  wire  Randomizer_33_clock; // @[GameLogic.scala 130:24]
  wire  Randomizer_33_reset; // @[GameLogic.scala 130:24]
  wire [1:0] Randomizer_33_io_out; // @[GameLogic.scala 130:24]
  wire  Randomizer_34_clock; // @[GameLogic.scala 107:24]
  wire  Randomizer_34_reset; // @[GameLogic.scala 107:24]
  wire [9:0] Randomizer_34_io_out; // @[GameLogic.scala 107:24]
  wire  Randomizer_35_clock; // @[GameLogic.scala 108:25]
  wire  Randomizer_35_reset; // @[GameLogic.scala 108:25]
  wire [5:0] Randomizer_35_io_out; // @[GameLogic.scala 108:25]
  wire  Randomizer_36_clock; // @[GameLogic.scala 107:24]
  wire  Randomizer_36_reset; // @[GameLogic.scala 107:24]
  wire [9:0] Randomizer_36_io_out; // @[GameLogic.scala 107:24]
  wire  Randomizer_37_clock; // @[GameLogic.scala 108:25]
  wire  Randomizer_37_reset; // @[GameLogic.scala 108:25]
  wire [5:0] Randomizer_37_io_out; // @[GameLogic.scala 108:25]
  wire  Randomizer_38_clock; // @[GameLogic.scala 107:24]
  wire  Randomizer_38_reset; // @[GameLogic.scala 107:24]
  wire [9:0] Randomizer_38_io_out; // @[GameLogic.scala 107:24]
  wire  Randomizer_39_clock; // @[GameLogic.scala 108:25]
  wire  Randomizer_39_reset; // @[GameLogic.scala 108:25]
  wire [5:0] Randomizer_39_io_out; // @[GameLogic.scala 108:25]
  wire  Randomizer_40_clock; // @[GameLogic.scala 130:24]
  wire  Randomizer_40_reset; // @[GameLogic.scala 130:24]
  wire [1:0] Randomizer_40_io_out; // @[GameLogic.scala 130:24]
  wire  Randomizer_41_clock; // @[GameLogic.scala 107:24]
  wire  Randomizer_41_reset; // @[GameLogic.scala 107:24]
  wire [9:0] Randomizer_41_io_out; // @[GameLogic.scala 107:24]
  wire  Randomizer_42_clock; // @[GameLogic.scala 108:25]
  wire  Randomizer_42_reset; // @[GameLogic.scala 108:25]
  wire [5:0] Randomizer_42_io_out; // @[GameLogic.scala 108:25]
  wire  Randomizer_43_clock; // @[GameLogic.scala 107:24]
  wire  Randomizer_43_reset; // @[GameLogic.scala 107:24]
  wire [9:0] Randomizer_43_io_out; // @[GameLogic.scala 107:24]
  wire  Randomizer_44_clock; // @[GameLogic.scala 108:25]
  wire  Randomizer_44_reset; // @[GameLogic.scala 108:25]
  wire [5:0] Randomizer_44_io_out; // @[GameLogic.scala 108:25]
  wire  Randomizer_45_clock; // @[GameLogic.scala 107:24]
  wire  Randomizer_45_reset; // @[GameLogic.scala 107:24]
  wire [9:0] Randomizer_45_io_out; // @[GameLogic.scala 107:24]
  wire  Randomizer_46_clock; // @[GameLogic.scala 108:25]
  wire  Randomizer_46_reset; // @[GameLogic.scala 108:25]
  wire [5:0] Randomizer_46_io_out; // @[GameLogic.scala 108:25]
  reg  planetUp; // @[GameLogic.scala 359:25]
  reg [10:0] Xstart_0; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_1; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_2; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_3; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_4; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_5; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_6; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_7; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_8; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_9; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_10; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_11; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_12; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_13; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_14; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_15; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_16; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_17; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_18; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_19; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_20; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_21; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_22; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_23; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_24; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_25; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_26; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_27; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_28; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_29; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_30; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_31; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_32; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_33; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_41; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_42; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_43; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_44; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_45; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_46; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_47; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_48; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_49; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_50; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_51; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_122; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_123; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_124; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_125; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_126; // @[GameLogic.scala 424:23]
  reg [10:0] Xstart_127; // @[GameLogic.scala 424:23]
  reg [10:0] Ystart_0; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_1; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_2; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_3; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_4; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_5; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_6; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_7; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_8; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_9; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_10; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_11; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_12; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_13; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_14; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_15; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_16; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_17; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_18; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_19; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_20; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_21; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_22; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_23; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_24; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_25; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_26; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_27; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_28; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_29; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_30; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_31; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_32; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_33; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_41; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_42; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_43; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_122; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_123; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_124; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_125; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_126; // @[GameLogic.scala 509:23]
  reg [10:0] Ystart_127; // @[GameLogic.scala 509:23]
  reg  spriteVisibleReg_0; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_1; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_2; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_3; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_4; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_5; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_6; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_7; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_8; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_9; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_10; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_11; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_12; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_13; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_14; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_15; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_16; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_17; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_18; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_19; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_20; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_21; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_22; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_23; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_24; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_25; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_26; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_27; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_28; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_29; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_30; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_31; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_32; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_33; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_41; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_42; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_43; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_44; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_45; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_46; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_47; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_48; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_49; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_50; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_51; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_55; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_56; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_57; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_61; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_62; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_63; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_64; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_65; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_66; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_70; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_71; // @[GameLogic.scala 620:33]
  reg  spriteVisibleReg_72; // @[GameLogic.scala 620:33]
  reg  spriteFlipVerticalReg_122; // @[GameLogic.scala 622:38]
  reg  spriteFlipVerticalReg_123; // @[GameLogic.scala 622:38]
  reg  spriteFlipVerticalReg_124; // @[GameLogic.scala 622:38]
  reg  spriteFlipVerticalReg_125; // @[GameLogic.scala 622:38]
  reg  spriteFlipVerticalReg_126; // @[GameLogic.scala 622:38]
  reg  spriteFlipVerticalReg_127; // @[GameLogic.scala 622:38]
  reg  btnCReg; // @[GameLogic.scala 623:24]
  reg [9:0] viewX; // @[GameLogic.scala 648:22]
  reg [3:0] stateReg; // @[GameLogic.scala 667:25]
  reg [9:0] shotCnt; // @[GameLogic.scala 670:24]
  reg  shotLoad; // @[GameLogic.scala 671:25]
  reg [2:0] shotCntBig; // @[GameLogic.scala 672:27]
  reg [2:0] shotCntFast; // @[GameLogic.scala 673:28]
  reg  shotPop_0; // @[GameLogic.scala 674:24]
  reg  shotPop_1; // @[GameLogic.scala 674:24]
  reg  shotPop_2; // @[GameLogic.scala 674:24]
  reg  shotPop_3; // @[GameLogic.scala 674:24]
  reg  shotPop_4; // @[GameLogic.scala 674:24]
  reg  shotInteract_0; // @[GameLogic.scala 675:29]
  reg  shotInteract_1; // @[GameLogic.scala 675:29]
  reg  shotInteract_2; // @[GameLogic.scala 675:29]
  reg  shotInteract_3; // @[GameLogic.scala 675:29]
  reg  shotInteract_4; // @[GameLogic.scala 675:29]
  reg  astInteract_0; // @[GameLogic.scala 676:28]
  reg  astInteract_1; // @[GameLogic.scala 676:28]
  reg  astInteract_2; // @[GameLogic.scala 676:28]
  reg  astInteract_3; // @[GameLogic.scala 676:28]
  reg  astInteract_4; // @[GameLogic.scala 676:28]
  reg  astInteract_5; // @[GameLogic.scala 676:28]
  reg  astInteract_6; // @[GameLogic.scala 676:28]
  reg  astInteract_7; // @[GameLogic.scala 676:28]
  reg  astInteract_8; // @[GameLogic.scala 676:28]
  reg  astInteract_9; // @[GameLogic.scala 676:28]
  reg  astInteract_10; // @[GameLogic.scala 676:28]
  reg  shipInteract; // @[GameLogic.scala 677:29]
  reg  die_0; // @[GameLogic.scala 679:20]
  reg  die_1; // @[GameLogic.scala 679:20]
  reg  die_2; // @[GameLogic.scala 679:20]
  reg  die_3; // @[GameLogic.scala 679:20]
  reg  die_4; // @[GameLogic.scala 679:20]
  reg  die_5; // @[GameLogic.scala 679:20]
  reg  die_6; // @[GameLogic.scala 679:20]
  reg  die_7; // @[GameLogic.scala 679:20]
  reg  die_8; // @[GameLogic.scala 679:20]
  reg  die_9; // @[GameLogic.scala 679:20]
  reg  die_10; // @[GameLogic.scala 679:20]
  reg  kill_0_0; // @[GameLogic.scala 680:21]
  reg  kill_0_1; // @[GameLogic.scala 680:21]
  reg  kill_0_2; // @[GameLogic.scala 680:21]
  reg  kill_0_3; // @[GameLogic.scala 680:21]
  reg  kill_0_4; // @[GameLogic.scala 680:21]
  reg  kill_1_0; // @[GameLogic.scala 680:21]
  reg  kill_1_1; // @[GameLogic.scala 680:21]
  reg  kill_1_2; // @[GameLogic.scala 680:21]
  reg  kill_1_3; // @[GameLogic.scala 680:21]
  reg  kill_1_4; // @[GameLogic.scala 680:21]
  reg  kill_2_0; // @[GameLogic.scala 680:21]
  reg  kill_2_1; // @[GameLogic.scala 680:21]
  reg  kill_2_2; // @[GameLogic.scala 680:21]
  reg  kill_2_3; // @[GameLogic.scala 680:21]
  reg  kill_2_4; // @[GameLogic.scala 680:21]
  reg  kill_3_0; // @[GameLogic.scala 680:21]
  reg  kill_3_1; // @[GameLogic.scala 680:21]
  reg  kill_3_2; // @[GameLogic.scala 680:21]
  reg  kill_3_3; // @[GameLogic.scala 680:21]
  reg  kill_3_4; // @[GameLogic.scala 680:21]
  reg  kill_4_0; // @[GameLogic.scala 680:21]
  reg  kill_4_1; // @[GameLogic.scala 680:21]
  reg  kill_4_2; // @[GameLogic.scala 680:21]
  reg  kill_4_3; // @[GameLogic.scala 680:21]
  reg  kill_4_4; // @[GameLogic.scala 680:21]
  reg  kill_5_0; // @[GameLogic.scala 680:21]
  reg  kill_5_1; // @[GameLogic.scala 680:21]
  reg  kill_5_2; // @[GameLogic.scala 680:21]
  reg  kill_5_3; // @[GameLogic.scala 680:21]
  reg  kill_5_4; // @[GameLogic.scala 680:21]
  reg  kill_6_0; // @[GameLogic.scala 680:21]
  reg  kill_6_1; // @[GameLogic.scala 680:21]
  reg  kill_6_2; // @[GameLogic.scala 680:21]
  reg  kill_6_3; // @[GameLogic.scala 680:21]
  reg  kill_6_4; // @[GameLogic.scala 680:21]
  reg  kill_7_0; // @[GameLogic.scala 680:21]
  reg  kill_7_1; // @[GameLogic.scala 680:21]
  reg  kill_7_2; // @[GameLogic.scala 680:21]
  reg  kill_7_3; // @[GameLogic.scala 680:21]
  reg  kill_7_4; // @[GameLogic.scala 680:21]
  reg  kill_8_0; // @[GameLogic.scala 680:21]
  reg  kill_8_1; // @[GameLogic.scala 680:21]
  reg  kill_8_2; // @[GameLogic.scala 680:21]
  reg  kill_8_3; // @[GameLogic.scala 680:21]
  reg  kill_8_4; // @[GameLogic.scala 680:21]
  reg  kill_9_0; // @[GameLogic.scala 680:21]
  reg  kill_9_1; // @[GameLogic.scala 680:21]
  reg  kill_9_2; // @[GameLogic.scala 680:21]
  reg  kill_9_3; // @[GameLogic.scala 680:21]
  reg  kill_10_0; // @[GameLogic.scala 680:21]
  reg  kill_10_1; // @[GameLogic.scala 680:21]
  reg  kill_10_2; // @[GameLogic.scala 680:21]
  reg  kill_10_3; // @[GameLogic.scala 680:21]
  reg  kill_10_4; // @[GameLogic.scala 680:21]
  reg [3:0] hp; // @[GameLogic.scala 682:19]
  reg [4:0] planetHp; // @[GameLogic.scala 683:25]
  reg [5:0] spwnProt; // @[GameLogic.scala 684:25]
  reg  show; // @[GameLogic.scala 685:21]
  reg  blink; // @[GameLogic.scala 686:22]
  reg [7:0] secCnt; // @[GameLogic.scala 687:23]
  reg [2:0] level; // @[GameLogic.scala 688:22]
  reg  start; // @[GameLogic.scala 689:22]
  reg  levelCng; // @[GameLogic.scala 690:25]
  reg [3:0] cngCnt; // @[GameLogic.scala 691:23]
  reg [9:0] cnt; // @[GameLogic.scala 693:20]
  wire  _T_25 = $signed(cnt) == 10'sh1d; // @[GameLogic.scala 694:17]
  wire  _T_26 = $signed(cnt) == 10'sh3b; // @[GameLogic.scala 694:33]
  wire  cng = _T_25 | _T_26; // @[GameLogic.scala 694:26]
  reg [6:0] count1; // @[GameLogic.scala 698:23]
  reg [6:0] count3; // @[GameLogic.scala 700:23]
  reg [7:0] count4; // @[GameLogic.scala 701:23]
  reg [7:0] count5; // @[GameLogic.scala 702:23]
  wire  _T_27 = ~show; // @[GameLogic.scala 706:26]
  wire  _T_28 = ~shipInteract; // @[GameLogic.scala 708:8]
  wire  _T_29 = _T_28 & blink; // @[GameLogic.scala 708:22]
  wire  _GEN_0 = _T_29 ? 1'h0 : show; // @[GameLogic.scala 708:32]
  wire  _GEN_1 = _T_29 ? 1'h0 : _T_27; // @[GameLogic.scala 708:32]
  wire [8:0] _T_33 = 8'sh0 / 8'sh2; // @[GameLogic.scala 714:66]
  wire [10:0] _GEN_4379 = {{2{_T_33[8]}},_T_33}; // @[GameLogic.scala 714:51]
  wire [10:0] _T_43 = $signed(Ystart_0) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_71 = $signed(Ystart_2) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_85 = $signed(Ystart_3) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_99 = $signed(Ystart_4) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_113 = $signed(Ystart_5) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_127 = $signed(Ystart_6) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [7:0] _T_130 = 8'sh20 - 8'sh8; // @[GameLogic.scala 714:57]
  wire [8:0] _T_131 = $signed(_T_130) / 8'sh2; // @[GameLogic.scala 714:66]
  wire [10:0] _GEN_4393 = {{2{_T_131[8]}},_T_131}; // @[GameLogic.scala 714:51]
  wire [10:0] _T_141 = $signed(Ystart_7) + $signed(_GEN_4393); // @[GameLogic.scala 715:51]
  wire [7:0] _T_144 = 8'sh20 - 8'sh10; // @[GameLogic.scala 714:57]
  wire [8:0] _T_145 = $signed(_T_144) / 8'sh2; // @[GameLogic.scala 714:66]
  wire [10:0] _GEN_4395 = {{2{_T_145[8]}},_T_145}; // @[GameLogic.scala 714:51]
  wire [10:0] _T_155 = $signed(Ystart_8) + $signed(_GEN_4395); // @[GameLogic.scala 715:51]
  wire [7:0] _T_158 = 8'sh20 - 8'sh1c; // @[GameLogic.scala 714:57]
  wire [8:0] _T_159 = $signed(_T_158) / 8'sh2; // @[GameLogic.scala 714:66]
  wire [10:0] _GEN_4397 = {{2{_T_159[8]}},_T_159}; // @[GameLogic.scala 714:51]
  wire [10:0] _T_169 = $signed(Ystart_9) + $signed(_GEN_4397); // @[GameLogic.scala 715:51]
  wire [10:0] _T_183 = $signed(Ystart_10) + $signed(_GEN_4397); // @[GameLogic.scala 715:51]
  wire [10:0] _T_197 = $signed(Ystart_11) + $signed(_GEN_4397); // @[GameLogic.scala 715:51]
  wire [10:0] _T_211 = $signed(Ystart_12) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_225 = $signed(Ystart_13) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_239 = $signed(Ystart_14) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_253 = $signed(Ystart_15) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [10:0] _T_267 = $signed(Ystart_16) + $signed(_GEN_4379); // @[GameLogic.scala 715:51]
  wire [7:0] _T_270 = 8'sh20 - 8'sh60; // @[GameLogic.scala 714:57]
  wire [8:0] _T_271 = $signed(_T_270) / 8'sh2; // @[GameLogic.scala 714:66]
  wire [10:0] _GEN_4413 = {{2{_T_271[8]}},_T_271}; // @[GameLogic.scala 714:51]
  wire [10:0] _T_281 = $signed(Ystart_17) + $signed(_GEN_4413); // @[GameLogic.scala 715:51]
  wire  _T_282 = hp <= 4'h0; // @[GameLogic.scala 342:13]
  wire  _T_283 = cngCnt == 4'h0; // @[GameLogic.scala 345:40]
  wire  _T_284 = cngCnt == 4'h1; // @[GameLogic.scala 346:40]
  wire  _T_285 = cngCnt == 4'h2; // @[GameLogic.scala 347:40]
  wire  _GEN_4 = _T_282 & _T_283; // @[GameLogic.scala 342:21]
  wire  _GEN_5 = _T_282 & _T_284; // @[GameLogic.scala 342:21]
  wire  _GEN_6 = _T_282 & _T_285; // @[GameLogic.scala 342:21]
  wire [11:0] _T_287 = {{1{Xstart_17[10]}},Xstart_17}; // @[GameLogic.scala 410:44]
  wire [10:0] _T_289 = _T_287[10:0]; // @[GameLogic.scala 410:44]
  wire [11:0] _T_290 = {{1{Ystart_17[10]}},Ystart_17}; // @[GameLogic.scala 411:44]
  wire [10:0] _T_292 = _T_290[10:0]; // @[GameLogic.scala 411:44]
  wire [10:0] _T_295 = $signed(Xstart_17) + 11'sh20; // @[GameLogic.scala 410:44]
  wire [10:0] _T_301 = $signed(Xstart_17) + 11'sh40; // @[GameLogic.scala 410:44]
  wire [10:0] _T_310 = $signed(Ystart_17) + 11'sh20; // @[GameLogic.scala 411:44]
  wire [10:0] _T_328 = $signed(Ystart_17) + 11'sh40; // @[GameLogic.scala 411:44]
  wire  _T_341 = planetHp < 5'h1; // @[GameLogic.scala 417:19]
  wire  _GEN_8 = _T_341 ? 1'h0 : astInteract_0; // @[GameLogic.scala 417:26]
  wire  _GEN_9 = _T_341 ? 1'h0 : spriteVisibleReg_7; // @[GameLogic.scala 417:26]
  wire  _GEN_10 = _T_341 ? 1'h0 : astInteract_1; // @[GameLogic.scala 417:26]
  wire  _GEN_11 = _T_341 ? 1'h0 : spriteVisibleReg_8; // @[GameLogic.scala 417:26]
  wire  _GEN_12 = _T_341 ? 1'h0 : astInteract_2; // @[GameLogic.scala 417:26]
  wire  _GEN_13 = _T_341 ? 1'h0 : spriteVisibleReg_9; // @[GameLogic.scala 417:26]
  wire  _GEN_14 = _T_341 ? 1'h0 : astInteract_3; // @[GameLogic.scala 417:26]
  wire  _GEN_15 = _T_341 ? 1'h0 : spriteVisibleReg_10; // @[GameLogic.scala 417:26]
  wire  _GEN_16 = _T_341 ? 1'h0 : astInteract_4; // @[GameLogic.scala 417:26]
  wire  _GEN_17 = _T_341 ? 1'h0 : spriteVisibleReg_11; // @[GameLogic.scala 417:26]
  wire  _GEN_18 = _T_341 ? 1'h0 : astInteract_5; // @[GameLogic.scala 417:26]
  wire  _GEN_19 = _T_341 ? 1'h0 : spriteVisibleReg_12; // @[GameLogic.scala 417:26]
  wire  _GEN_20 = _T_341 ? 1'h0 : astInteract_6; // @[GameLogic.scala 417:26]
  wire  _GEN_21 = _T_341 ? 1'h0 : spriteVisibleReg_13; // @[GameLogic.scala 417:26]
  wire  _GEN_22 = _T_341 ? 1'h0 : astInteract_7; // @[GameLogic.scala 417:26]
  wire  _GEN_23 = _T_341 ? 1'h0 : spriteVisibleReg_14; // @[GameLogic.scala 417:26]
  wire  _GEN_24 = _T_341 ? 1'h0 : astInteract_8; // @[GameLogic.scala 417:26]
  wire  _GEN_25 = _T_341 ? 1'h0 : spriteVisibleReg_15; // @[GameLogic.scala 417:26]
  wire  _GEN_26 = _T_341 ? 1'h0 : astInteract_9; // @[GameLogic.scala 417:26]
  wire  _GEN_27 = _T_341 ? 1'h0 : spriteVisibleReg_16; // @[GameLogic.scala 417:26]
  wire  _GEN_28 = _T_341 ? 1'h0 : astInteract_10; // @[GameLogic.scala 417:26]
  wire  _GEN_29 = _T_341 ? 1'h0 : spriteVisibleReg_17; // @[GameLogic.scala 417:26]
  wire  _T_342 = 4'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_343 = 4'h1 == stateReg; // @[Conditional.scala 37:30]
  wire [9:0] _T_346 = viewX + 10'h2; // @[GameLogic.scala 733:22]
  wire [10:0] _T_349 = $signed(Xstart_2) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_352 = $signed(Xstart_3) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_355 = $signed(Xstart_4) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_358 = $signed(Xstart_5) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_361 = $signed(Xstart_6) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_364 = $signed(Xstart_7) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_367 = $signed(Xstart_8) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_370 = $signed(Xstart_9) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_373 = $signed(Xstart_10) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_376 = $signed(Xstart_11) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_379 = $signed(Xstart_12) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_382 = $signed(Xstart_13) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_385 = $signed(Xstart_14) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_388 = $signed(Xstart_15) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_391 = $signed(Xstart_16) - 11'sh2; // @[GameLogic.scala 742:40]
  wire [10:0] _T_394 = $signed(Xstart_17) - 11'sh2; // @[GameLogic.scala 742:40]
  wire  _T_396 = viewX >= 10'h20; // @[GameLogic.scala 746:18]
  wire [9:0] _T_399 = viewX - 10'h20; // @[GameLogic.scala 748:24]
  wire [9:0] _T_402 = _T_399 + 10'h2; // @[GameLogic.scala 748:43]
  wire [6:0] _T_404 = count1 + 7'h1; // @[GameLogic.scala 752:28]
  wire  _T_405 = 4'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_406 = count1 >= 7'h1a; // @[GameLogic.scala 760:19]
  wire  _T_407 = viewX >= 10'h16; // @[GameLogic.scala 765:18]
  wire  _T_408 = count4 == 8'h1; // @[GameLogic.scala 767:21]
  wire  _T_409 = count3 < 7'h9; // @[GameLogic.scala 768:23]
  wire [2:0] _T_411 = level - 3'h1; // @[GameLogic.scala 769:53]
  wire [5:0] _T_412 = _T_411 * 3'h5; // @[GameLogic.scala 769:60]
  wire [5:0] _T_414 = 6'hc + _T_412; // @[GameLogic.scala 769:44]
  wire [7:0] _GEN_4415 = {{1'd0}, count1}; // @[GameLogic.scala 770:48]
  wire [7:0] _T_416 = 8'h8f - _GEN_4415; // @[GameLogic.scala 770:48]
  wire [12:0] _T_417 = count3 * 7'h28; // @[GameLogic.scala 770:66]
  wire [12:0] _GEN_4416 = {{5'd0}, _T_416}; // @[GameLogic.scala 770:57]
  wire [12:0] _T_419 = _GEN_4416 + _T_417; // @[GameLogic.scala 770:57]
  wire [6:0] _T_421 = count3 + 7'h1; // @[GameLogic.scala 773:30]
  wire [5:0] _GEN_37 = _T_409 ? _T_414 : 6'h0; // @[GameLogic.scala 768:30]
  wire [12:0] _GEN_38 = _T_409 ? _T_419 : 13'h0; // @[GameLogic.scala 768:30]
  wire [6:0] _GEN_40 = _T_409 ? _T_421 : 7'h0; // @[GameLogic.scala 768:30]
  wire [5:0] _GEN_42 = _T_408 ? _GEN_37 : 6'h0; // @[GameLogic.scala 767:30]
  wire [12:0] _GEN_43 = _T_408 ? _GEN_38 : 13'h0; // @[GameLogic.scala 767:30]
  wire  _GEN_44 = _T_408 & _T_409; // @[GameLogic.scala 767:30]
  wire [5:0] _GEN_47 = _T_407 ? _GEN_42 : 6'h0; // @[GameLogic.scala 765:27]
  wire [12:0] _GEN_48 = _T_407 ? _GEN_43 : 13'h0; // @[GameLogic.scala 765:27]
  wire  _GEN_49 = _T_407 & _GEN_44; // @[GameLogic.scala 765:27]
  wire  _T_422 = viewX < 10'h16; // @[GameLogic.scala 782:19]
  wire  _T_423 = viewX >= 10'hb; // @[GameLogic.scala 782:37]
  wire  _T_424 = _T_422 & _T_423; // @[GameLogic.scala 782:27]
  wire [5:0] _T_430 = 6'hb + _T_412; // @[GameLogic.scala 785:42]
  wire [5:0] _GEN_52 = _T_409 ? _T_430 : _GEN_47; // @[GameLogic.scala 784:28]
  wire [12:0] _GEN_53 = _T_409 ? _T_419 : _GEN_48; // @[GameLogic.scala 784:28]
  wire  _GEN_54 = _T_409 | _GEN_49; // @[GameLogic.scala 784:28]
  wire [5:0] _GEN_57 = _T_424 ? _GEN_52 : _GEN_47; // @[GameLogic.scala 782:47]
  wire [12:0] _GEN_58 = _T_424 ? _GEN_53 : _GEN_48; // @[GameLogic.scala 782:47]
  wire  _GEN_59 = _T_424 ? _GEN_54 : _GEN_49; // @[GameLogic.scala 782:47]
  wire  _T_438 = viewX < 10'hb; // @[GameLogic.scala 796:18]
  wire [5:0] _T_444 = 6'ha + _T_412; // @[GameLogic.scala 799:42]
  wire [5:0] _GEN_62 = _T_409 ? _T_444 : _GEN_57; // @[GameLogic.scala 798:28]
  wire [12:0] _GEN_63 = _T_409 ? _T_419 : _GEN_58; // @[GameLogic.scala 798:28]
  wire  _GEN_64 = _T_409 | _GEN_59; // @[GameLogic.scala 798:28]
  wire [5:0] _GEN_67 = _T_438 ? _GEN_62 : _GEN_57; // @[GameLogic.scala 796:26]
  wire [12:0] _GEN_68 = _T_438 ? _GEN_63 : _GEN_58; // @[GameLogic.scala 796:26]
  wire  _GEN_69 = _T_438 ? _GEN_64 : _GEN_59; // @[GameLogic.scala 796:26]
  wire  _T_452 = 4'h3 == stateReg; // @[Conditional.scala 37:30]
  wire [5:0] _T_465 = 6'he + _T_412; // @[GameLogic.scala 821:42]
  wire [7:0] _T_467 = 8'h90 - _GEN_4415; // @[GameLogic.scala 822:46]
  wire [12:0] _GEN_4422 = {{5'd0}, _T_467}; // @[GameLogic.scala 822:55]
  wire [12:0] _T_470 = _GEN_4422 + _T_417; // @[GameLogic.scala 822:55]
  wire [5:0] _GEN_76 = _T_409 ? _T_465 : 6'h0; // @[GameLogic.scala 820:28]
  wire [12:0] _GEN_77 = _T_409 ? _T_470 : 13'h0; // @[GameLogic.scala 820:28]
  wire [5:0] _GEN_82 = _T_424 ? _GEN_76 : 6'h0; // @[GameLogic.scala 819:47]
  wire [12:0] _GEN_83 = _T_424 ? _GEN_77 : 13'h0; // @[GameLogic.scala 819:47]
  wire  _GEN_84 = _T_424 & _T_409; // @[GameLogic.scala 819:47]
  wire [5:0] _T_479 = 6'hd + _T_412; // @[GameLogic.scala 834:42]
  wire [5:0] _GEN_88 = _T_409 ? _T_479 : _GEN_82; // @[GameLogic.scala 833:28]
  wire [12:0] _GEN_89 = _T_409 ? _T_470 : _GEN_83; // @[GameLogic.scala 833:28]
  wire  _GEN_90 = _T_409 | _GEN_84; // @[GameLogic.scala 833:28]
  wire [5:0] _GEN_93 = _T_438 ? _GEN_88 : _GEN_82; // @[GameLogic.scala 832:26]
  wire [12:0] _GEN_94 = _T_438 ? _GEN_89 : _GEN_83; // @[GameLogic.scala 832:26]
  wire  _GEN_95 = _T_438 ? _GEN_90 : _GEN_84; // @[GameLogic.scala 832:26]
  wire  _T_487 = 4'h4 == stateReg; // @[Conditional.scala 37:30]
  wire [7:0] _T_495 = 8'h91 - _GEN_4415; // @[GameLogic.scala 849:44]
  wire [12:0] _GEN_4426 = {{5'd0}, _T_495}; // @[GameLogic.scala 849:53]
  wire [12:0] _T_498 = _GEN_4426 + _T_417; // @[GameLogic.scala 849:53]
  wire  _T_501 = planetHp <= 5'h0; // @[GameLogic.scala 853:27]
  wire  _T_502 = level >= 3'h4; // @[GameLogic.scala 857:31]
  wire  _T_503 = $signed(secCnt) >= 8'sha; // @[GameLogic.scala 857:48]
  wire  _T_504 = _T_502 & _T_503; // @[GameLogic.scala 857:38]
  wire [12:0] _GEN_101 = _T_409 ? _T_498 : 13'h0; // @[GameLogic.scala 847:26]
  wire  _T_506 = 4'h5 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_507 = level < 3'h4; // @[GameLogic.scala 862:27]
  wire  _T_508 = start & _T_507; // @[GameLogic.scala 862:18]
  wire [10:0] _T_511 = $signed(Xstart_7) - 11'sh4; // @[GameLogic.scala 306:44]
  wire  _T_512 = planetHp >= 5'h1; // @[GameLogic.scala 307:19]
  wire  _T_513 = $signed(Xstart_7) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_514 = $signed(secCnt) >= 8'sh5; // @[GameLogic.scala 203:45]
  wire  _T_515 = _T_513 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4427 = {{4{Randomizer_1_io_out[6]}},Randomizer_1_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_522 = $signed(_GEN_4427) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire [9:0] _T_523 = viewX; // @[GameLogic.scala 210:47]
  wire [10:0] _GEN_4428 = {{1{_T_523[9]}},_T_523}; // @[GameLogic.scala 210:39]
  wire [10:0] _T_526 = 11'sh2c0 + $signed(_GEN_4428); // @[GameLogic.scala 210:39]
  wire [10:0] _GEN_105 = _T_502 ? $signed(_T_295) : $signed(_T_526); // @[GameLogic.scala 206:26]
  wire  _GEN_107 = _T_515 | _GEN_8; // @[GameLogic.scala 203:53]
  wire  _GEN_108 = _T_515 | _GEN_9; // @[GameLogic.scala 203:53]
  wire  _GEN_115 = kill_0_3 & shotInteract_0; // @[GameLogic.scala 169:41]
  wire  _GEN_116 = kill_0_3 ? shotPop_0 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_117 = kill_0_3 & spriteVisibleReg_2; // @[GameLogic.scala 169:41]
  wire  _GEN_119 = kill_0_0 ? _GEN_115 : shotInteract_0; // @[GameLogic.scala 167:39]
  wire  _GEN_120 = kill_0_0 ? _GEN_116 : shotPop_0; // @[GameLogic.scala 167:39]
  wire  _GEN_121 = kill_0_0 ? _GEN_117 : spriteVisibleReg_2; // @[GameLogic.scala 167:39]
  wire  _GEN_123 = kill_0_3 & shotInteract_1; // @[GameLogic.scala 169:41]
  wire  _GEN_124 = kill_0_3 ? shotPop_1 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_125 = kill_0_3 & spriteVisibleReg_3; // @[GameLogic.scala 169:41]
  wire  _GEN_127 = kill_0_1 ? _GEN_123 : shotInteract_1; // @[GameLogic.scala 167:39]
  wire  _GEN_128 = kill_0_1 ? _GEN_124 : shotPop_1; // @[GameLogic.scala 167:39]
  wire  _GEN_129 = kill_0_1 ? _GEN_125 : spriteVisibleReg_3; // @[GameLogic.scala 167:39]
  wire  _GEN_131 = kill_0_3 & shotInteract_2; // @[GameLogic.scala 169:41]
  wire  _GEN_132 = kill_0_3 ? shotPop_2 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_133 = kill_0_3 & spriteVisibleReg_4; // @[GameLogic.scala 169:41]
  wire  _GEN_135 = kill_0_2 ? _GEN_131 : shotInteract_2; // @[GameLogic.scala 167:39]
  wire  _GEN_136 = kill_0_2 ? _GEN_132 : shotPop_2; // @[GameLogic.scala 167:39]
  wire  _GEN_137 = kill_0_2 ? _GEN_133 : spriteVisibleReg_4; // @[GameLogic.scala 167:39]
  wire  _GEN_139 = kill_0_3 & shotInteract_3; // @[GameLogic.scala 169:41]
  wire  _GEN_140 = kill_0_3 ? shotPop_3 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_141 = kill_0_3 & spriteVisibleReg_5; // @[GameLogic.scala 169:41]
  wire  _GEN_143 = kill_0_3 ? _GEN_139 : shotInteract_3; // @[GameLogic.scala 167:39]
  wire  _GEN_144 = kill_0_3 ? _GEN_140 : shotPop_3; // @[GameLogic.scala 167:39]
  wire  _GEN_145 = kill_0_3 ? _GEN_141 : spriteVisibleReg_5; // @[GameLogic.scala 167:39]
  wire  _GEN_147 = kill_0_3 & shotInteract_4; // @[GameLogic.scala 169:41]
  wire  _GEN_148 = kill_0_3 ? shotPop_4 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_149 = kill_0_3 & spriteVisibleReg_6; // @[GameLogic.scala 169:41]
  wire  _GEN_151 = kill_0_4 ? _GEN_147 : shotInteract_4; // @[GameLogic.scala 167:39]
  wire  _GEN_152 = kill_0_4 ? _GEN_148 : shotPop_4; // @[GameLogic.scala 167:39]
  wire  _GEN_153 = kill_0_4 ? _GEN_149 : spriteVisibleReg_6; // @[GameLogic.scala 167:39]
  wire [10:0] _T_529 = $signed(Xstart_8) - 11'sh4; // @[GameLogic.scala 306:44]
  wire  _T_531 = $signed(Xstart_8) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_533 = _T_531 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4429 = {{4{Randomizer_3_io_out[6]}},Randomizer_3_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_540 = $signed(_GEN_4429) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_157 = _T_533 | _GEN_10; // @[GameLogic.scala 203:53]
  wire  _GEN_158 = _T_533 | _GEN_11; // @[GameLogic.scala 203:53]
  wire  _GEN_165 = kill_1_3 & _GEN_119; // @[GameLogic.scala 169:41]
  wire  _GEN_166 = kill_1_3 ? _GEN_120 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_167 = kill_1_3 & _GEN_121; // @[GameLogic.scala 169:41]
  wire  _GEN_169 = kill_1_0 ? _GEN_165 : _GEN_119; // @[GameLogic.scala 167:39]
  wire  _GEN_170 = kill_1_0 ? _GEN_166 : _GEN_120; // @[GameLogic.scala 167:39]
  wire  _GEN_171 = kill_1_0 ? _GEN_167 : _GEN_121; // @[GameLogic.scala 167:39]
  wire  _GEN_173 = kill_1_3 & _GEN_127; // @[GameLogic.scala 169:41]
  wire  _GEN_174 = kill_1_3 ? _GEN_128 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_175 = kill_1_3 & _GEN_129; // @[GameLogic.scala 169:41]
  wire  _GEN_177 = kill_1_1 ? _GEN_173 : _GEN_127; // @[GameLogic.scala 167:39]
  wire  _GEN_178 = kill_1_1 ? _GEN_174 : _GEN_128; // @[GameLogic.scala 167:39]
  wire  _GEN_179 = kill_1_1 ? _GEN_175 : _GEN_129; // @[GameLogic.scala 167:39]
  wire  _GEN_181 = kill_1_3 & _GEN_135; // @[GameLogic.scala 169:41]
  wire  _GEN_182 = kill_1_3 ? _GEN_136 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_183 = kill_1_3 & _GEN_137; // @[GameLogic.scala 169:41]
  wire  _GEN_185 = kill_1_2 ? _GEN_181 : _GEN_135; // @[GameLogic.scala 167:39]
  wire  _GEN_186 = kill_1_2 ? _GEN_182 : _GEN_136; // @[GameLogic.scala 167:39]
  wire  _GEN_187 = kill_1_2 ? _GEN_183 : _GEN_137; // @[GameLogic.scala 167:39]
  wire  _GEN_189 = kill_1_3 & _GEN_143; // @[GameLogic.scala 169:41]
  wire  _GEN_190 = kill_1_3 ? _GEN_144 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_191 = kill_1_3 & _GEN_145; // @[GameLogic.scala 169:41]
  wire  _GEN_193 = kill_1_3 ? _GEN_189 : _GEN_143; // @[GameLogic.scala 167:39]
  wire  _GEN_194 = kill_1_3 ? _GEN_190 : _GEN_144; // @[GameLogic.scala 167:39]
  wire  _GEN_195 = kill_1_3 ? _GEN_191 : _GEN_145; // @[GameLogic.scala 167:39]
  wire  _GEN_197 = kill_1_3 & _GEN_151; // @[GameLogic.scala 169:41]
  wire  _GEN_198 = kill_1_3 ? _GEN_152 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_199 = kill_1_3 & _GEN_153; // @[GameLogic.scala 169:41]
  wire  _GEN_201 = kill_1_4 ? _GEN_197 : _GEN_151; // @[GameLogic.scala 167:39]
  wire  _GEN_202 = kill_1_4 ? _GEN_198 : _GEN_152; // @[GameLogic.scala 167:39]
  wire  _GEN_203 = kill_1_4 ? _GEN_199 : _GEN_153; // @[GameLogic.scala 167:39]
  wire [10:0] _T_547 = $signed(Xstart_9) - 11'sh4; // @[GameLogic.scala 306:44]
  wire  _T_549 = $signed(Xstart_9) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_551 = _T_549 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4431 = {{4{Randomizer_5_io_out[6]}},Randomizer_5_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_558 = $signed(_GEN_4431) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_207 = _T_551 | _GEN_12; // @[GameLogic.scala 203:53]
  wire  _GEN_208 = _T_551 | _GEN_13; // @[GameLogic.scala 203:53]
  wire  _GEN_215 = kill_2_3 & _GEN_169; // @[GameLogic.scala 169:41]
  wire  _GEN_216 = kill_2_3 ? _GEN_170 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_217 = kill_2_3 & _GEN_171; // @[GameLogic.scala 169:41]
  wire  _GEN_219 = kill_2_0 ? _GEN_215 : _GEN_169; // @[GameLogic.scala 167:39]
  wire  _GEN_220 = kill_2_0 ? _GEN_216 : _GEN_170; // @[GameLogic.scala 167:39]
  wire  _GEN_221 = kill_2_0 ? _GEN_217 : _GEN_171; // @[GameLogic.scala 167:39]
  wire  _GEN_223 = kill_2_3 & _GEN_177; // @[GameLogic.scala 169:41]
  wire  _GEN_224 = kill_2_3 ? _GEN_178 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_225 = kill_2_3 & _GEN_179; // @[GameLogic.scala 169:41]
  wire  _GEN_227 = kill_2_1 ? _GEN_223 : _GEN_177; // @[GameLogic.scala 167:39]
  wire  _GEN_228 = kill_2_1 ? _GEN_224 : _GEN_178; // @[GameLogic.scala 167:39]
  wire  _GEN_229 = kill_2_1 ? _GEN_225 : _GEN_179; // @[GameLogic.scala 167:39]
  wire  _GEN_231 = kill_2_3 & _GEN_185; // @[GameLogic.scala 169:41]
  wire  _GEN_232 = kill_2_3 ? _GEN_186 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_233 = kill_2_3 & _GEN_187; // @[GameLogic.scala 169:41]
  wire  _GEN_235 = kill_2_2 ? _GEN_231 : _GEN_185; // @[GameLogic.scala 167:39]
  wire  _GEN_236 = kill_2_2 ? _GEN_232 : _GEN_186; // @[GameLogic.scala 167:39]
  wire  _GEN_237 = kill_2_2 ? _GEN_233 : _GEN_187; // @[GameLogic.scala 167:39]
  wire  _GEN_239 = kill_2_3 & _GEN_193; // @[GameLogic.scala 169:41]
  wire  _GEN_240 = kill_2_3 ? _GEN_194 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_241 = kill_2_3 & _GEN_195; // @[GameLogic.scala 169:41]
  wire  _GEN_243 = kill_2_3 ? _GEN_239 : _GEN_193; // @[GameLogic.scala 167:39]
  wire  _GEN_244 = kill_2_3 ? _GEN_240 : _GEN_194; // @[GameLogic.scala 167:39]
  wire  _GEN_245 = kill_2_3 ? _GEN_241 : _GEN_195; // @[GameLogic.scala 167:39]
  wire  _GEN_247 = kill_2_3 & _GEN_201; // @[GameLogic.scala 169:41]
  wire  _GEN_248 = kill_2_3 ? _GEN_202 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_249 = kill_2_3 & _GEN_203; // @[GameLogic.scala 169:41]
  wire  _GEN_251 = kill_2_4 ? _GEN_247 : _GEN_201; // @[GameLogic.scala 167:39]
  wire  _GEN_252 = kill_2_4 ? _GEN_248 : _GEN_202; // @[GameLogic.scala 167:39]
  wire  _GEN_253 = kill_2_4 ? _GEN_249 : _GEN_203; // @[GameLogic.scala 167:39]
  wire  _T_563 = level >= 3'h1; // @[GameLogic.scala 866:31]
  wire  _T_566 = _T_502 & _T_514; // @[GameLogic.scala 866:56]
  wire  _GEN_259 = _T_508 ? _GEN_219 : shotInteract_0; // @[GameLogic.scala 862:34]
  wire  _GEN_260 = _T_508 ? _GEN_220 : shotPop_0; // @[GameLogic.scala 862:34]
  wire  _GEN_261 = _T_508 ? _GEN_221 : spriteVisibleReg_2; // @[GameLogic.scala 862:34]
  wire  _GEN_262 = _T_508 ? _GEN_227 : shotInteract_1; // @[GameLogic.scala 862:34]
  wire  _GEN_263 = _T_508 ? _GEN_228 : shotPop_1; // @[GameLogic.scala 862:34]
  wire  _GEN_264 = _T_508 ? _GEN_229 : spriteVisibleReg_3; // @[GameLogic.scala 862:34]
  wire  _GEN_265 = _T_508 ? _GEN_235 : shotInteract_2; // @[GameLogic.scala 862:34]
  wire  _GEN_266 = _T_508 ? _GEN_236 : shotPop_2; // @[GameLogic.scala 862:34]
  wire  _GEN_267 = _T_508 ? _GEN_237 : spriteVisibleReg_4; // @[GameLogic.scala 862:34]
  wire  _GEN_268 = _T_508 ? _GEN_243 : shotInteract_3; // @[GameLogic.scala 862:34]
  wire  _GEN_269 = _T_508 ? _GEN_244 : shotPop_3; // @[GameLogic.scala 862:34]
  wire  _GEN_270 = _T_508 ? _GEN_245 : spriteVisibleReg_5; // @[GameLogic.scala 862:34]
  wire  _GEN_271 = _T_508 ? _GEN_251 : shotInteract_4; // @[GameLogic.scala 862:34]
  wire  _GEN_272 = _T_508 ? _GEN_252 : shotPop_4; // @[GameLogic.scala 862:34]
  wire  _GEN_273 = _T_508 ? _GEN_253 : spriteVisibleReg_6; // @[GameLogic.scala 862:34]
  wire  _T_571 = 4'h6 == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_574 = $signed(Xstart_10) - 11'sh4; // @[GameLogic.scala 306:44]
  wire  _T_576 = $signed(Xstart_10) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_578 = _T_576 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4433 = {{4{Randomizer_7_io_out[6]}},Randomizer_7_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_585 = $signed(_GEN_4433) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_285 = _T_578 | _GEN_14; // @[GameLogic.scala 203:53]
  wire  _GEN_286 = _T_578 | _GEN_15; // @[GameLogic.scala 203:53]
  wire  _GEN_293 = kill_3_3 & shotInteract_0; // @[GameLogic.scala 169:41]
  wire  _GEN_294 = kill_3_3 ? shotPop_0 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_295 = kill_3_3 & spriteVisibleReg_2; // @[GameLogic.scala 169:41]
  wire  _GEN_297 = kill_3_0 ? _GEN_293 : shotInteract_0; // @[GameLogic.scala 167:39]
  wire  _GEN_298 = kill_3_0 ? _GEN_294 : shotPop_0; // @[GameLogic.scala 167:39]
  wire  _GEN_299 = kill_3_0 ? _GEN_295 : spriteVisibleReg_2; // @[GameLogic.scala 167:39]
  wire  _GEN_301 = kill_3_3 & shotInteract_1; // @[GameLogic.scala 169:41]
  wire  _GEN_302 = kill_3_3 ? shotPop_1 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_303 = kill_3_3 & spriteVisibleReg_3; // @[GameLogic.scala 169:41]
  wire  _GEN_305 = kill_3_1 ? _GEN_301 : shotInteract_1; // @[GameLogic.scala 167:39]
  wire  _GEN_306 = kill_3_1 ? _GEN_302 : shotPop_1; // @[GameLogic.scala 167:39]
  wire  _GEN_307 = kill_3_1 ? _GEN_303 : spriteVisibleReg_3; // @[GameLogic.scala 167:39]
  wire  _GEN_309 = kill_3_3 & shotInteract_2; // @[GameLogic.scala 169:41]
  wire  _GEN_310 = kill_3_3 ? shotPop_2 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_311 = kill_3_3 & spriteVisibleReg_4; // @[GameLogic.scala 169:41]
  wire  _GEN_313 = kill_3_2 ? _GEN_309 : shotInteract_2; // @[GameLogic.scala 167:39]
  wire  _GEN_314 = kill_3_2 ? _GEN_310 : shotPop_2; // @[GameLogic.scala 167:39]
  wire  _GEN_315 = kill_3_2 ? _GEN_311 : spriteVisibleReg_4; // @[GameLogic.scala 167:39]
  wire  _GEN_317 = kill_3_3 & shotInteract_3; // @[GameLogic.scala 169:41]
  wire  _GEN_318 = kill_3_3 ? shotPop_3 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_319 = kill_3_3 & spriteVisibleReg_5; // @[GameLogic.scala 169:41]
  wire  _GEN_321 = kill_3_3 ? _GEN_317 : shotInteract_3; // @[GameLogic.scala 167:39]
  wire  _GEN_322 = kill_3_3 ? _GEN_318 : shotPop_3; // @[GameLogic.scala 167:39]
  wire  _GEN_323 = kill_3_3 ? _GEN_319 : spriteVisibleReg_5; // @[GameLogic.scala 167:39]
  wire  _GEN_325 = kill_3_3 & shotInteract_4; // @[GameLogic.scala 169:41]
  wire  _GEN_326 = kill_3_3 ? shotPop_4 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_327 = kill_3_3 & spriteVisibleReg_6; // @[GameLogic.scala 169:41]
  wire  _GEN_329 = kill_3_4 ? _GEN_325 : shotInteract_4; // @[GameLogic.scala 167:39]
  wire  _GEN_330 = kill_3_4 ? _GEN_326 : shotPop_4; // @[GameLogic.scala 167:39]
  wire  _GEN_331 = kill_3_4 ? _GEN_327 : spriteVisibleReg_6; // @[GameLogic.scala 167:39]
  wire [10:0] _T_592 = $signed(Xstart_11) - 11'sh5; // @[GameLogic.scala 306:44]
  wire  _T_594 = $signed(Xstart_11) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_596 = _T_594 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4435 = {{4{Randomizer_9_io_out[6]}},Randomizer_9_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_603 = $signed(_GEN_4435) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_335 = _T_596 | _GEN_16; // @[GameLogic.scala 203:53]
  wire  _GEN_336 = _T_596 | _GEN_17; // @[GameLogic.scala 203:53]
  wire  _GEN_343 = kill_4_3 & _GEN_297; // @[GameLogic.scala 169:41]
  wire  _GEN_344 = kill_4_3 ? _GEN_298 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_345 = kill_4_3 & _GEN_299; // @[GameLogic.scala 169:41]
  wire  _GEN_347 = kill_4_0 ? _GEN_343 : _GEN_297; // @[GameLogic.scala 167:39]
  wire  _GEN_348 = kill_4_0 ? _GEN_344 : _GEN_298; // @[GameLogic.scala 167:39]
  wire  _GEN_349 = kill_4_0 ? _GEN_345 : _GEN_299; // @[GameLogic.scala 167:39]
  wire  _GEN_351 = kill_4_3 & _GEN_305; // @[GameLogic.scala 169:41]
  wire  _GEN_352 = kill_4_3 ? _GEN_306 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_353 = kill_4_3 & _GEN_307; // @[GameLogic.scala 169:41]
  wire  _GEN_355 = kill_4_1 ? _GEN_351 : _GEN_305; // @[GameLogic.scala 167:39]
  wire  _GEN_356 = kill_4_1 ? _GEN_352 : _GEN_306; // @[GameLogic.scala 167:39]
  wire  _GEN_357 = kill_4_1 ? _GEN_353 : _GEN_307; // @[GameLogic.scala 167:39]
  wire  _GEN_359 = kill_4_3 & _GEN_313; // @[GameLogic.scala 169:41]
  wire  _GEN_360 = kill_4_3 ? _GEN_314 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_361 = kill_4_3 & _GEN_315; // @[GameLogic.scala 169:41]
  wire  _GEN_363 = kill_4_2 ? _GEN_359 : _GEN_313; // @[GameLogic.scala 167:39]
  wire  _GEN_364 = kill_4_2 ? _GEN_360 : _GEN_314; // @[GameLogic.scala 167:39]
  wire  _GEN_365 = kill_4_2 ? _GEN_361 : _GEN_315; // @[GameLogic.scala 167:39]
  wire  _GEN_367 = kill_4_3 & _GEN_321; // @[GameLogic.scala 169:41]
  wire  _GEN_368 = kill_4_3 ? _GEN_322 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_369 = kill_4_3 & _GEN_323; // @[GameLogic.scala 169:41]
  wire  _GEN_371 = kill_4_3 ? _GEN_367 : _GEN_321; // @[GameLogic.scala 167:39]
  wire  _GEN_372 = kill_4_3 ? _GEN_368 : _GEN_322; // @[GameLogic.scala 167:39]
  wire  _GEN_373 = kill_4_3 ? _GEN_369 : _GEN_323; // @[GameLogic.scala 167:39]
  wire  _GEN_375 = kill_4_3 & _GEN_329; // @[GameLogic.scala 169:41]
  wire  _GEN_376 = kill_4_3 ? _GEN_330 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_377 = kill_4_3 & _GEN_331; // @[GameLogic.scala 169:41]
  wire  _GEN_379 = kill_4_4 ? _GEN_375 : _GEN_329; // @[GameLogic.scala 167:39]
  wire  _GEN_380 = kill_4_4 ? _GEN_376 : _GEN_330; // @[GameLogic.scala 167:39]
  wire  _GEN_381 = kill_4_4 ? _GEN_377 : _GEN_331; // @[GameLogic.scala 167:39]
  wire [10:0] _T_610 = $signed(Xstart_12) - 11'sh5; // @[GameLogic.scala 306:44]
  wire  _T_612 = $signed(Xstart_12) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_614 = _T_612 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4437 = {{4{Randomizer_11_io_out[6]}},Randomizer_11_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_621 = $signed(_GEN_4437) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_385 = _T_614 | _GEN_18; // @[GameLogic.scala 203:53]
  wire  _GEN_386 = _T_614 | _GEN_19; // @[GameLogic.scala 203:53]
  wire  _GEN_393 = kill_5_3 & _GEN_347; // @[GameLogic.scala 169:41]
  wire  _GEN_394 = kill_5_3 ? _GEN_348 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_395 = kill_5_3 & _GEN_349; // @[GameLogic.scala 169:41]
  wire  _GEN_397 = kill_5_0 ? _GEN_393 : _GEN_347; // @[GameLogic.scala 167:39]
  wire  _GEN_398 = kill_5_0 ? _GEN_394 : _GEN_348; // @[GameLogic.scala 167:39]
  wire  _GEN_399 = kill_5_0 ? _GEN_395 : _GEN_349; // @[GameLogic.scala 167:39]
  wire  _GEN_401 = kill_5_3 & _GEN_355; // @[GameLogic.scala 169:41]
  wire  _GEN_402 = kill_5_3 ? _GEN_356 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_403 = kill_5_3 & _GEN_357; // @[GameLogic.scala 169:41]
  wire  _GEN_405 = kill_5_1 ? _GEN_401 : _GEN_355; // @[GameLogic.scala 167:39]
  wire  _GEN_406 = kill_5_1 ? _GEN_402 : _GEN_356; // @[GameLogic.scala 167:39]
  wire  _GEN_407 = kill_5_1 ? _GEN_403 : _GEN_357; // @[GameLogic.scala 167:39]
  wire  _GEN_409 = kill_5_3 & _GEN_363; // @[GameLogic.scala 169:41]
  wire  _GEN_410 = kill_5_3 ? _GEN_364 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_411 = kill_5_3 & _GEN_365; // @[GameLogic.scala 169:41]
  wire  _GEN_413 = kill_5_2 ? _GEN_409 : _GEN_363; // @[GameLogic.scala 167:39]
  wire  _GEN_414 = kill_5_2 ? _GEN_410 : _GEN_364; // @[GameLogic.scala 167:39]
  wire  _GEN_415 = kill_5_2 ? _GEN_411 : _GEN_365; // @[GameLogic.scala 167:39]
  wire  _GEN_417 = kill_5_3 & _GEN_371; // @[GameLogic.scala 169:41]
  wire  _GEN_418 = kill_5_3 ? _GEN_372 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_419 = kill_5_3 & _GEN_373; // @[GameLogic.scala 169:41]
  wire  _GEN_421 = kill_5_3 ? _GEN_417 : _GEN_371; // @[GameLogic.scala 167:39]
  wire  _GEN_422 = kill_5_3 ? _GEN_418 : _GEN_372; // @[GameLogic.scala 167:39]
  wire  _GEN_423 = kill_5_3 ? _GEN_419 : _GEN_373; // @[GameLogic.scala 167:39]
  wire  _GEN_425 = kill_5_3 & _GEN_379; // @[GameLogic.scala 169:41]
  wire  _GEN_426 = kill_5_3 ? _GEN_380 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_427 = kill_5_3 & _GEN_381; // @[GameLogic.scala 169:41]
  wire  _GEN_429 = kill_5_4 ? _GEN_425 : _GEN_379; // @[GameLogic.scala 167:39]
  wire  _GEN_430 = kill_5_4 ? _GEN_426 : _GEN_380; // @[GameLogic.scala 167:39]
  wire  _GEN_431 = kill_5_4 ? _GEN_427 : _GEN_381; // @[GameLogic.scala 167:39]
  wire  _T_626 = level >= 3'h2; // @[GameLogic.scala 877:29]
  wire  _T_628 = 4'h7 == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_631 = $signed(Xstart_13) - 11'sh5; // @[GameLogic.scala 306:44]
  wire  _T_633 = $signed(Xstart_13) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_635 = _T_633 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4439 = {{4{Randomizer_13_io_out[6]}},Randomizer_13_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_642 = $signed(_GEN_4439) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_435 = _T_635 | _GEN_20; // @[GameLogic.scala 203:53]
  wire  _GEN_436 = _T_635 | _GEN_21; // @[GameLogic.scala 203:53]
  wire  _GEN_443 = kill_6_3 & shotInteract_0; // @[GameLogic.scala 169:41]
  wire  _GEN_444 = kill_6_3 ? shotPop_0 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_445 = kill_6_3 & spriteVisibleReg_2; // @[GameLogic.scala 169:41]
  wire  _GEN_447 = kill_6_0 ? _GEN_443 : shotInteract_0; // @[GameLogic.scala 167:39]
  wire  _GEN_448 = kill_6_0 ? _GEN_444 : shotPop_0; // @[GameLogic.scala 167:39]
  wire  _GEN_449 = kill_6_0 ? _GEN_445 : spriteVisibleReg_2; // @[GameLogic.scala 167:39]
  wire  _GEN_451 = kill_6_3 & shotInteract_1; // @[GameLogic.scala 169:41]
  wire  _GEN_452 = kill_6_3 ? shotPop_1 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_453 = kill_6_3 & spriteVisibleReg_3; // @[GameLogic.scala 169:41]
  wire  _GEN_455 = kill_6_1 ? _GEN_451 : shotInteract_1; // @[GameLogic.scala 167:39]
  wire  _GEN_456 = kill_6_1 ? _GEN_452 : shotPop_1; // @[GameLogic.scala 167:39]
  wire  _GEN_457 = kill_6_1 ? _GEN_453 : spriteVisibleReg_3; // @[GameLogic.scala 167:39]
  wire  _GEN_459 = kill_6_3 & shotInteract_2; // @[GameLogic.scala 169:41]
  wire  _GEN_460 = kill_6_3 ? shotPop_2 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_461 = kill_6_3 & spriteVisibleReg_4; // @[GameLogic.scala 169:41]
  wire  _GEN_463 = kill_6_2 ? _GEN_459 : shotInteract_2; // @[GameLogic.scala 167:39]
  wire  _GEN_464 = kill_6_2 ? _GEN_460 : shotPop_2; // @[GameLogic.scala 167:39]
  wire  _GEN_465 = kill_6_2 ? _GEN_461 : spriteVisibleReg_4; // @[GameLogic.scala 167:39]
  wire  _GEN_467 = kill_6_3 & shotInteract_3; // @[GameLogic.scala 169:41]
  wire  _GEN_468 = kill_6_3 ? shotPop_3 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_469 = kill_6_3 & spriteVisibleReg_5; // @[GameLogic.scala 169:41]
  wire  _GEN_471 = kill_6_3 ? _GEN_467 : shotInteract_3; // @[GameLogic.scala 167:39]
  wire  _GEN_472 = kill_6_3 ? _GEN_468 : shotPop_3; // @[GameLogic.scala 167:39]
  wire  _GEN_473 = kill_6_3 ? _GEN_469 : spriteVisibleReg_5; // @[GameLogic.scala 167:39]
  wire  _GEN_475 = kill_6_3 & shotInteract_4; // @[GameLogic.scala 169:41]
  wire  _GEN_476 = kill_6_3 ? shotPop_4 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_477 = kill_6_3 & spriteVisibleReg_6; // @[GameLogic.scala 169:41]
  wire  _GEN_479 = kill_6_4 ? _GEN_475 : shotInteract_4; // @[GameLogic.scala 167:39]
  wire  _GEN_480 = kill_6_4 ? _GEN_476 : shotPop_4; // @[GameLogic.scala 167:39]
  wire  _GEN_481 = kill_6_4 ? _GEN_477 : spriteVisibleReg_6; // @[GameLogic.scala 167:39]
  wire [10:0] _T_649 = $signed(Xstart_14) - 11'sh3; // @[GameLogic.scala 306:44]
  wire  _T_651 = $signed(Xstart_14) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_653 = _T_651 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4441 = {{4{Randomizer_15_io_out[6]}},Randomizer_15_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_660 = $signed(_GEN_4441) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_485 = _T_653 | _GEN_22; // @[GameLogic.scala 203:53]
  wire  _GEN_486 = _T_653 | _GEN_23; // @[GameLogic.scala 203:53]
  wire  _GEN_493 = kill_7_3 & _GEN_447; // @[GameLogic.scala 169:41]
  wire  _GEN_494 = kill_7_3 ? _GEN_448 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_495 = kill_7_3 & _GEN_449; // @[GameLogic.scala 169:41]
  wire  _GEN_497 = kill_7_0 ? _GEN_493 : _GEN_447; // @[GameLogic.scala 167:39]
  wire  _GEN_498 = kill_7_0 ? _GEN_494 : _GEN_448; // @[GameLogic.scala 167:39]
  wire  _GEN_499 = kill_7_0 ? _GEN_495 : _GEN_449; // @[GameLogic.scala 167:39]
  wire  _GEN_501 = kill_7_3 & _GEN_455; // @[GameLogic.scala 169:41]
  wire  _GEN_502 = kill_7_3 ? _GEN_456 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_503 = kill_7_3 & _GEN_457; // @[GameLogic.scala 169:41]
  wire  _GEN_505 = kill_7_1 ? _GEN_501 : _GEN_455; // @[GameLogic.scala 167:39]
  wire  _GEN_506 = kill_7_1 ? _GEN_502 : _GEN_456; // @[GameLogic.scala 167:39]
  wire  _GEN_507 = kill_7_1 ? _GEN_503 : _GEN_457; // @[GameLogic.scala 167:39]
  wire  _GEN_509 = kill_7_3 & _GEN_463; // @[GameLogic.scala 169:41]
  wire  _GEN_510 = kill_7_3 ? _GEN_464 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_511 = kill_7_3 & _GEN_465; // @[GameLogic.scala 169:41]
  wire  _GEN_513 = kill_7_2 ? _GEN_509 : _GEN_463; // @[GameLogic.scala 167:39]
  wire  _GEN_514 = kill_7_2 ? _GEN_510 : _GEN_464; // @[GameLogic.scala 167:39]
  wire  _GEN_515 = kill_7_2 ? _GEN_511 : _GEN_465; // @[GameLogic.scala 167:39]
  wire  _GEN_517 = kill_7_3 & _GEN_471; // @[GameLogic.scala 169:41]
  wire  _GEN_518 = kill_7_3 ? _GEN_472 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_519 = kill_7_3 & _GEN_473; // @[GameLogic.scala 169:41]
  wire  _GEN_521 = kill_7_3 ? _GEN_517 : _GEN_471; // @[GameLogic.scala 167:39]
  wire  _GEN_522 = kill_7_3 ? _GEN_518 : _GEN_472; // @[GameLogic.scala 167:39]
  wire  _GEN_523 = kill_7_3 ? _GEN_519 : _GEN_473; // @[GameLogic.scala 167:39]
  wire  _GEN_525 = kill_7_3 & _GEN_479; // @[GameLogic.scala 169:41]
  wire  _GEN_526 = kill_7_3 ? _GEN_480 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_527 = kill_7_3 & _GEN_481; // @[GameLogic.scala 169:41]
  wire  _GEN_529 = kill_7_4 ? _GEN_525 : _GEN_479; // @[GameLogic.scala 167:39]
  wire  _GEN_530 = kill_7_4 ? _GEN_526 : _GEN_480; // @[GameLogic.scala 167:39]
  wire  _GEN_531 = kill_7_4 ? _GEN_527 : _GEN_481; // @[GameLogic.scala 167:39]
  wire [10:0] _T_667 = $signed(Xstart_15) - 11'sh3; // @[GameLogic.scala 306:44]
  wire  _T_669 = $signed(Xstart_15) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_671 = _T_669 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4443 = {{4{Randomizer_17_io_out[6]}},Randomizer_17_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_678 = $signed(_GEN_4443) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_535 = _T_671 | _GEN_24; // @[GameLogic.scala 203:53]
  wire  _GEN_536 = _T_671 | _GEN_25; // @[GameLogic.scala 203:53]
  wire  _GEN_543 = kill_8_3 & _GEN_497; // @[GameLogic.scala 169:41]
  wire  _GEN_544 = kill_8_3 ? _GEN_498 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_545 = kill_8_3 & _GEN_499; // @[GameLogic.scala 169:41]
  wire  _GEN_547 = kill_8_0 ? _GEN_543 : _GEN_497; // @[GameLogic.scala 167:39]
  wire  _GEN_548 = kill_8_0 ? _GEN_544 : _GEN_498; // @[GameLogic.scala 167:39]
  wire  _GEN_549 = kill_8_0 ? _GEN_545 : _GEN_499; // @[GameLogic.scala 167:39]
  wire  _GEN_551 = kill_8_3 & _GEN_505; // @[GameLogic.scala 169:41]
  wire  _GEN_552 = kill_8_3 ? _GEN_506 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_553 = kill_8_3 & _GEN_507; // @[GameLogic.scala 169:41]
  wire  _GEN_555 = kill_8_1 ? _GEN_551 : _GEN_505; // @[GameLogic.scala 167:39]
  wire  _GEN_556 = kill_8_1 ? _GEN_552 : _GEN_506; // @[GameLogic.scala 167:39]
  wire  _GEN_557 = kill_8_1 ? _GEN_553 : _GEN_507; // @[GameLogic.scala 167:39]
  wire  _GEN_559 = kill_8_3 & _GEN_513; // @[GameLogic.scala 169:41]
  wire  _GEN_560 = kill_8_3 ? _GEN_514 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_561 = kill_8_3 & _GEN_515; // @[GameLogic.scala 169:41]
  wire  _GEN_563 = kill_8_2 ? _GEN_559 : _GEN_513; // @[GameLogic.scala 167:39]
  wire  _GEN_564 = kill_8_2 ? _GEN_560 : _GEN_514; // @[GameLogic.scala 167:39]
  wire  _GEN_565 = kill_8_2 ? _GEN_561 : _GEN_515; // @[GameLogic.scala 167:39]
  wire  _GEN_567 = kill_8_3 & _GEN_521; // @[GameLogic.scala 169:41]
  wire  _GEN_568 = kill_8_3 ? _GEN_522 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_569 = kill_8_3 & _GEN_523; // @[GameLogic.scala 169:41]
  wire  _GEN_571 = kill_8_3 ? _GEN_567 : _GEN_521; // @[GameLogic.scala 167:39]
  wire  _GEN_572 = kill_8_3 ? _GEN_568 : _GEN_522; // @[GameLogic.scala 167:39]
  wire  _GEN_573 = kill_8_3 ? _GEN_569 : _GEN_523; // @[GameLogic.scala 167:39]
  wire  _GEN_575 = kill_8_3 & _GEN_529; // @[GameLogic.scala 169:41]
  wire  _GEN_576 = kill_8_3 ? _GEN_530 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_577 = kill_8_3 & _GEN_531; // @[GameLogic.scala 169:41]
  wire  _GEN_579 = kill_8_4 ? _GEN_575 : _GEN_529; // @[GameLogic.scala 167:39]
  wire  _GEN_580 = kill_8_4 ? _GEN_576 : _GEN_530; // @[GameLogic.scala 167:39]
  wire  _GEN_581 = kill_8_4 ? _GEN_577 : _GEN_531; // @[GameLogic.scala 167:39]
  wire  _T_683 = level >= 3'h3; // @[GameLogic.scala 884:29]
  wire  _T_685 = 4'h8 == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_688 = $signed(Xstart_16) - 11'sh4; // @[GameLogic.scala 181:44]
  wire  _T_689 = planetHp > 5'h0; // @[GameLogic.scala 182:19]
  wire  _T_690 = $signed(Xstart_16) <= 11'sh2; // @[GameLogic.scala 203:28]
  wire  _T_692 = _T_690 & _T_514; // @[GameLogic.scala 203:35]
  wire [10:0] _GEN_4445 = {{4{Randomizer_19_io_out[6]}},Randomizer_19_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_699 = $signed(_GEN_4445) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_585 = _T_692 | _GEN_26; // @[GameLogic.scala 203:53]
  wire  _GEN_586 = _T_692 | _GEN_27; // @[GameLogic.scala 203:53]
  wire  _GEN_593 = kill_9_0 ? 1'h0 : shotInteract_0; // @[GameLogic.scala 186:39]
  wire  _GEN_594 = kill_9_0 | shotPop_0; // @[GameLogic.scala 186:39]
  wire  _GEN_595 = kill_9_0 ? 1'h0 : spriteVisibleReg_2; // @[GameLogic.scala 186:39]
  wire  _GEN_596 = kill_9_1 ? 1'h0 : shotInteract_1; // @[GameLogic.scala 186:39]
  wire  _GEN_597 = kill_9_1 | shotPop_1; // @[GameLogic.scala 186:39]
  wire  _GEN_598 = kill_9_1 ? 1'h0 : spriteVisibleReg_3; // @[GameLogic.scala 186:39]
  wire  _GEN_599 = kill_9_2 ? 1'h0 : shotInteract_2; // @[GameLogic.scala 186:39]
  wire  _GEN_600 = kill_9_2 | shotPop_2; // @[GameLogic.scala 186:39]
  wire  _GEN_601 = kill_9_2 ? 1'h0 : spriteVisibleReg_4; // @[GameLogic.scala 186:39]
  wire  _T_706 = 4'h9 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_707 = $signed(secCnt) >= 8'shb; // @[GameLogic.scala 893:19]
  wire [10:0] _GEN_4447 = {{4{Randomizer_21_io_out[6]}},Randomizer_21_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_721 = $signed(_GEN_4447) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire [10:0] _GEN_4449 = {{4{Randomizer_23_io_out[6]}},Randomizer_23_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_739 = $signed(_GEN_4449) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire [10:0] _GEN_4451 = {{4{Randomizer_25_io_out[6]}},Randomizer_25_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_757 = $signed(_GEN_4451) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire [10:0] _GEN_4453 = {{4{Randomizer_27_io_out[6]}},Randomizer_27_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_775 = $signed(_GEN_4453) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_674 = kill_4_3 & _GEN_219; // @[GameLogic.scala 169:41]
  wire  _GEN_675 = kill_4_3 ? _GEN_220 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_676 = kill_4_3 & _GEN_221; // @[GameLogic.scala 169:41]
  wire  _GEN_678 = kill_4_0 ? _GEN_674 : _GEN_219; // @[GameLogic.scala 167:39]
  wire  _GEN_679 = kill_4_0 ? _GEN_675 : _GEN_220; // @[GameLogic.scala 167:39]
  wire  _GEN_680 = kill_4_0 ? _GEN_676 : _GEN_221; // @[GameLogic.scala 167:39]
  wire  _GEN_682 = kill_4_3 & _GEN_227; // @[GameLogic.scala 169:41]
  wire  _GEN_683 = kill_4_3 ? _GEN_228 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_684 = kill_4_3 & _GEN_229; // @[GameLogic.scala 169:41]
  wire  _GEN_686 = kill_4_1 ? _GEN_682 : _GEN_227; // @[GameLogic.scala 167:39]
  wire  _GEN_687 = kill_4_1 ? _GEN_683 : _GEN_228; // @[GameLogic.scala 167:39]
  wire  _GEN_688 = kill_4_1 ? _GEN_684 : _GEN_229; // @[GameLogic.scala 167:39]
  wire  _GEN_690 = kill_4_3 & _GEN_235; // @[GameLogic.scala 169:41]
  wire  _GEN_691 = kill_4_3 ? _GEN_236 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_692 = kill_4_3 & _GEN_237; // @[GameLogic.scala 169:41]
  wire  _GEN_694 = kill_4_2 ? _GEN_690 : _GEN_235; // @[GameLogic.scala 167:39]
  wire  _GEN_695 = kill_4_2 ? _GEN_691 : _GEN_236; // @[GameLogic.scala 167:39]
  wire  _GEN_696 = kill_4_2 ? _GEN_692 : _GEN_237; // @[GameLogic.scala 167:39]
  wire  _GEN_698 = kill_4_3 & _GEN_243; // @[GameLogic.scala 169:41]
  wire  _GEN_699 = kill_4_3 ? _GEN_244 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_700 = kill_4_3 & _GEN_245; // @[GameLogic.scala 169:41]
  wire  _GEN_702 = kill_4_3 ? _GEN_698 : _GEN_243; // @[GameLogic.scala 167:39]
  wire  _GEN_703 = kill_4_3 ? _GEN_699 : _GEN_244; // @[GameLogic.scala 167:39]
  wire  _GEN_704 = kill_4_3 ? _GEN_700 : _GEN_245; // @[GameLogic.scala 167:39]
  wire  _GEN_706 = kill_4_3 & _GEN_251; // @[GameLogic.scala 169:41]
  wire  _GEN_707 = kill_4_3 ? _GEN_252 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_708 = kill_4_3 & _GEN_253; // @[GameLogic.scala 169:41]
  wire  _GEN_710 = kill_4_4 ? _GEN_706 : _GEN_251; // @[GameLogic.scala 167:39]
  wire  _GEN_711 = kill_4_4 ? _GEN_707 : _GEN_252; // @[GameLogic.scala 167:39]
  wire  _GEN_712 = kill_4_4 ? _GEN_708 : _GEN_253; // @[GameLogic.scala 167:39]
  wire [10:0] _GEN_4455 = {{4{Randomizer_29_io_out[6]}},Randomizer_29_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_793 = $signed(_GEN_4455) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_724 = kill_5_3 & _GEN_678; // @[GameLogic.scala 169:41]
  wire  _GEN_725 = kill_5_3 ? _GEN_679 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_726 = kill_5_3 & _GEN_680; // @[GameLogic.scala 169:41]
  wire  _GEN_728 = kill_5_0 ? _GEN_724 : _GEN_678; // @[GameLogic.scala 167:39]
  wire  _GEN_729 = kill_5_0 ? _GEN_725 : _GEN_679; // @[GameLogic.scala 167:39]
  wire  _GEN_730 = kill_5_0 ? _GEN_726 : _GEN_680; // @[GameLogic.scala 167:39]
  wire  _GEN_732 = kill_5_3 & _GEN_686; // @[GameLogic.scala 169:41]
  wire  _GEN_733 = kill_5_3 ? _GEN_687 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_734 = kill_5_3 & _GEN_688; // @[GameLogic.scala 169:41]
  wire  _GEN_736 = kill_5_1 ? _GEN_732 : _GEN_686; // @[GameLogic.scala 167:39]
  wire  _GEN_737 = kill_5_1 ? _GEN_733 : _GEN_687; // @[GameLogic.scala 167:39]
  wire  _GEN_738 = kill_5_1 ? _GEN_734 : _GEN_688; // @[GameLogic.scala 167:39]
  wire  _GEN_740 = kill_5_3 & _GEN_694; // @[GameLogic.scala 169:41]
  wire  _GEN_741 = kill_5_3 ? _GEN_695 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_742 = kill_5_3 & _GEN_696; // @[GameLogic.scala 169:41]
  wire  _GEN_744 = kill_5_2 ? _GEN_740 : _GEN_694; // @[GameLogic.scala 167:39]
  wire  _GEN_745 = kill_5_2 ? _GEN_741 : _GEN_695; // @[GameLogic.scala 167:39]
  wire  _GEN_746 = kill_5_2 ? _GEN_742 : _GEN_696; // @[GameLogic.scala 167:39]
  wire  _GEN_748 = kill_5_3 & _GEN_702; // @[GameLogic.scala 169:41]
  wire  _GEN_749 = kill_5_3 ? _GEN_703 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_750 = kill_5_3 & _GEN_704; // @[GameLogic.scala 169:41]
  wire  _GEN_752 = kill_5_3 ? _GEN_748 : _GEN_702; // @[GameLogic.scala 167:39]
  wire  _GEN_753 = kill_5_3 ? _GEN_749 : _GEN_703; // @[GameLogic.scala 167:39]
  wire  _GEN_754 = kill_5_3 ? _GEN_750 : _GEN_704; // @[GameLogic.scala 167:39]
  wire  _GEN_756 = kill_5_3 & _GEN_710; // @[GameLogic.scala 169:41]
  wire  _GEN_757 = kill_5_3 ? _GEN_711 : 1'h1; // @[GameLogic.scala 169:41]
  wire  _GEN_758 = kill_5_3 & _GEN_712; // @[GameLogic.scala 169:41]
  wire  _GEN_760 = kill_5_4 ? _GEN_756 : _GEN_710; // @[GameLogic.scala 167:39]
  wire  _GEN_761 = kill_5_4 ? _GEN_757 : _GEN_711; // @[GameLogic.scala 167:39]
  wire  _GEN_762 = kill_5_4 ? _GEN_758 : _GEN_712; // @[GameLogic.scala 167:39]
  wire [10:0] _GEN_4457 = {{4{Randomizer_31_io_out[6]}},Randomizer_31_io_out}; // @[GameLogic.scala 208:51]
  wire [10:0] _T_811 = $signed(_GEN_4457) + $signed(Ystart_17); // @[GameLogic.scala 208:51]
  wire  _GEN_774 = kill_9_0 ? 1'h0 : _GEN_728; // @[GameLogic.scala 186:39]
  wire  _GEN_775 = kill_9_0 | _GEN_729; // @[GameLogic.scala 186:39]
  wire  _GEN_776 = kill_9_0 ? 1'h0 : _GEN_730; // @[GameLogic.scala 186:39]
  wire  _GEN_777 = kill_9_1 ? 1'h0 : _GEN_736; // @[GameLogic.scala 186:39]
  wire  _GEN_778 = kill_9_1 | _GEN_737; // @[GameLogic.scala 186:39]
  wire  _GEN_779 = kill_9_1 ? 1'h0 : _GEN_738; // @[GameLogic.scala 186:39]
  wire  _GEN_780 = kill_9_2 ? 1'h0 : _GEN_744; // @[GameLogic.scala 186:39]
  wire  _GEN_781 = kill_9_2 | _GEN_745; // @[GameLogic.scala 186:39]
  wire  _GEN_782 = kill_9_2 ? 1'h0 : _GEN_746; // @[GameLogic.scala 186:39]
  wire  _GEN_789 = _T_707 ? _GEN_774 : shotInteract_0; // @[GameLogic.scala 893:27]
  wire  _GEN_790 = _T_707 ? _GEN_775 : shotPop_0; // @[GameLogic.scala 893:27]
  wire  _GEN_791 = _T_707 ? _GEN_776 : spriteVisibleReg_2; // @[GameLogic.scala 893:27]
  wire  _GEN_792 = _T_707 ? _GEN_777 : shotInteract_1; // @[GameLogic.scala 893:27]
  wire  _GEN_793 = _T_707 ? _GEN_778 : shotPop_1; // @[GameLogic.scala 893:27]
  wire  _GEN_794 = _T_707 ? _GEN_779 : spriteVisibleReg_3; // @[GameLogic.scala 893:27]
  wire  _GEN_795 = _T_707 ? _GEN_780 : shotInteract_2; // @[GameLogic.scala 893:27]
  wire  _GEN_796 = _T_707 ? _GEN_781 : shotPop_2; // @[GameLogic.scala 893:27]
  wire  _GEN_797 = _T_707 ? _GEN_782 : spriteVisibleReg_4; // @[GameLogic.scala 893:27]
  wire  _GEN_798 = _T_707 ? _GEN_752 : shotInteract_3; // @[GameLogic.scala 893:27]
  wire  _GEN_799 = _T_707 ? _GEN_753 : shotPop_3; // @[GameLogic.scala 893:27]
  wire  _GEN_800 = _T_707 ? _GEN_754 : spriteVisibleReg_5; // @[GameLogic.scala 893:27]
  wire  _GEN_801 = _T_707 ? _GEN_760 : shotInteract_4; // @[GameLogic.scala 893:27]
  wire  _GEN_802 = _T_707 ? _GEN_761 : shotPop_4; // @[GameLogic.scala 893:27]
  wire  _GEN_803 = _T_707 ? _GEN_762 : spriteVisibleReg_6; // @[GameLogic.scala 893:27]
  wire  _T_816 = $signed(Ystart_17) <= 11'sh60; // @[GameLogic.scala 362:25]
  wire  _T_817 = $signed(Ystart_17) >= 11'sh120; // @[GameLogic.scala 364:31]
  wire  _GEN_824 = _T_817 | planetUp; // @[GameLogic.scala 364:43]
  wire  _GEN_825 = _T_816 ? 1'h0 : _GEN_824; // @[GameLogic.scala 362:37]
  wire  _T_818 = ~planetUp; // @[GameLogic.scala 367:44]
  wire [4:0] _T_821 = 5'sh0 - 5'sh1; // @[GameLogic.scala 367:69]
  wire [4:0] _T_822 = _T_818 ? $signed(5'sh1) : $signed(_T_821); // @[GameLogic.scala 367:43]
  wire [10:0] _GEN_4459 = {{6{_T_822[4]}},_T_822}; // @[GameLogic.scala 367:38]
  wire [10:0] _T_825 = $signed(Ystart_17) + $signed(_GEN_4459); // @[GameLogic.scala 367:38]
  wire  _T_826 = $signed(Xstart_17) > 11'sh1e0; // @[GameLogic.scala 368:42]
  wire [10:0] _T_829 = $signed(Xstart_17) - 11'sh1; // @[GameLogic.scala 368:69]
  wire  _T_831 = ~astInteract_10; // @[GameLogic.scala 375:10]
  wire  _T_834 = _T_514 & _T_689; // @[GameLogic.scala 376:26]
  wire [9:0] _T_841 = 10'sh160 - 10'sh40; // @[GameLogic.scala 380:54]
  wire  _T_842 = $signed(Randomizer_32_io_out) >= $signed(_T_841); // @[GameLogic.scala 380:45]
  wire [9:0] _T_846 = _T_842 ? $signed(_T_841) : $signed(Randomizer_32_io_out); // @[GameLogic.scala 380:30]
  wire  _GEN_826 = _T_834 | _GEN_28; // @[GameLogic.scala 376:45]
  wire  _GEN_827 = _T_834 | _GEN_29; // @[GameLogic.scala 376:45]
  wire [4:0] _T_849 = planetHp - 5'h1; // @[GameLogic.scala 390:32]
  wire [4:0] _GEN_834 = _T_689 ? _T_849 : planetHp; // @[GameLogic.scala 389:30]
  wire [4:0] _GEN_835 = kill_10_0 ? _GEN_834 : planetHp; // @[GameLogic.scala 387:36]
  wire  _GEN_836 = kill_10_0 ? 1'h0 : _GEN_789; // @[GameLogic.scala 387:36]
  wire  _GEN_837 = kill_10_0 | _GEN_790; // @[GameLogic.scala 387:36]
  wire  _GEN_838 = kill_10_0 ? 1'h0 : _GEN_791; // @[GameLogic.scala 387:36]
  wire [4:0] _GEN_839 = _T_689 ? _T_849 : _GEN_835; // @[GameLogic.scala 389:30]
  wire [4:0] _GEN_840 = kill_10_1 ? _GEN_839 : _GEN_835; // @[GameLogic.scala 387:36]
  wire  _GEN_841 = kill_10_1 ? 1'h0 : _GEN_792; // @[GameLogic.scala 387:36]
  wire  _GEN_842 = kill_10_1 | _GEN_793; // @[GameLogic.scala 387:36]
  wire  _GEN_843 = kill_10_1 ? 1'h0 : _GEN_794; // @[GameLogic.scala 387:36]
  wire  _GEN_846 = kill_10_2 ? 1'h0 : _GEN_795; // @[GameLogic.scala 387:36]
  wire  _GEN_847 = kill_10_2 | _GEN_796; // @[GameLogic.scala 387:36]
  wire  _GEN_848 = kill_10_2 ? 1'h0 : _GEN_797; // @[GameLogic.scala 387:36]
  wire  _GEN_851 = kill_10_3 ? 1'h0 : _GEN_798; // @[GameLogic.scala 387:36]
  wire  _GEN_852 = kill_10_3 | _GEN_799; // @[GameLogic.scala 387:36]
  wire  _GEN_853 = kill_10_3 ? 1'h0 : _GEN_800; // @[GameLogic.scala 387:36]
  wire  _GEN_856 = kill_10_4 ? 1'h0 : _GEN_801; // @[GameLogic.scala 387:36]
  wire  _GEN_857 = kill_10_4 | _GEN_802; // @[GameLogic.scala 387:36]
  wire  _GEN_858 = kill_10_4 ? 1'h0 : _GEN_803; // @[GameLogic.scala 387:36]
  wire  _T_863 = 4'ha == stateReg; // @[Conditional.scala 37:30]
  wire  _T_864 = hp > 4'h0; // @[GameLogic.scala 911:15]
  wire  _T_865 = $signed(Ystart_0) < 11'sh160; // @[GameLogic.scala 914:30]
  wire [10:0] _T_868 = $signed(Ystart_0) + 11'sh3; // @[GameLogic.scala 915:44]
  wire  _T_869 = $signed(Ystart_0) > 11'sh60; // @[GameLogic.scala 919:32]
  wire [10:0] _T_872 = $signed(Ystart_0) - 11'sh3; // @[GameLogic.scala 920:46]
  wire [9:0] _T_875 = 10'sh1c0 - 10'sh10; // @[GameLogic.scala 924:42]
  wire [10:0] _GEN_4461 = {{1{_T_875[9]}},_T_875}; // @[GameLogic.scala 924:30]
  wire  _T_876 = $signed(Xstart_0) < $signed(_GEN_4461); // @[GameLogic.scala 924:30]
  wire [10:0] _T_879 = $signed(Xstart_0) + 11'sh3; // @[GameLogic.scala 925:44]
  wire  _T_883 = $signed(Xstart_0) > 11'sh21; // @[GameLogic.scala 930:32]
  wire [10:0] _T_886 = $signed(Xstart_0) - 11'sh3; // @[GameLogic.scala 931:46]
  wire  _T_887 = 4'hb == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_890 = $signed(Xstart_2) + 11'sha; // @[GameLogic.scala 942:64]
  wire  _T_891 = $signed(Xstart_2) >= 11'sh280; // @[GameLogic.scala 278:36]
  wire  _GEN_872 = _T_891 ? 1'h0 : spriteVisibleReg_2; // @[GameLogic.scala 278:49]
  wire  _GEN_873 = _T_891 ? 1'h0 : shotInteract_0; // @[GameLogic.scala 278:49]
  wire  _GEN_874 = _T_891 | shotPop_0; // @[GameLogic.scala 278:49]
  wire [10:0] _T_894 = $signed(Xstart_3) + 11'sha; // @[GameLogic.scala 942:64]
  wire  _T_895 = $signed(Xstart_3) >= 11'sh280; // @[GameLogic.scala 278:36]
  wire  _GEN_875 = _T_895 ? 1'h0 : spriteVisibleReg_3; // @[GameLogic.scala 278:49]
  wire  _GEN_876 = _T_895 ? 1'h0 : shotInteract_1; // @[GameLogic.scala 278:49]
  wire  _GEN_877 = _T_895 | shotPop_1; // @[GameLogic.scala 278:49]
  wire [10:0] _T_898 = $signed(Xstart_4) + 11'sha; // @[GameLogic.scala 942:64]
  wire  _T_899 = $signed(Xstart_4) >= 11'sh280; // @[GameLogic.scala 278:36]
  wire  _GEN_878 = _T_899 ? 1'h0 : spriteVisibleReg_4; // @[GameLogic.scala 278:49]
  wire  _GEN_879 = _T_899 ? 1'h0 : shotInteract_2; // @[GameLogic.scala 278:49]
  wire  _GEN_880 = _T_899 | shotPop_2; // @[GameLogic.scala 278:49]
  wire [10:0] _T_902 = $signed(Xstart_5) + 11'sha; // @[GameLogic.scala 942:64]
  wire  _T_903 = $signed(Xstart_5) >= 11'sh280; // @[GameLogic.scala 278:36]
  wire  _GEN_881 = _T_903 ? 1'h0 : spriteVisibleReg_5; // @[GameLogic.scala 278:49]
  wire  _GEN_882 = _T_903 ? 1'h0 : shotInteract_3; // @[GameLogic.scala 278:49]
  wire  _GEN_883 = _T_903 | shotPop_3; // @[GameLogic.scala 278:49]
  wire [10:0] _T_906 = $signed(Xstart_6) + 11'sh1e; // @[GameLogic.scala 942:64]
  wire  _T_907 = $signed(Xstart_6) >= 11'sh280; // @[GameLogic.scala 278:36]
  wire  _GEN_884 = _T_907 ? 1'h0 : spriteVisibleReg_6; // @[GameLogic.scala 278:49]
  wire  _GEN_885 = _T_907 ? 1'h0 : shotInteract_4; // @[GameLogic.scala 278:49]
  wire  _GEN_886 = _T_907 | shotPop_4; // @[GameLogic.scala 278:49]
  wire  _T_909 = $signed(shotCntBig) > 3'sh0; // @[GameLogic.scala 946:37]
  wire  _T_910 = io_sw_1 & _T_909; // @[GameLogic.scala 946:23]
  wire  _T_912 = btnCReg & _T_909; // @[GameLogic.scala 258:18]
  wire  _GEN_887 = _T_912 | shotLoad; // @[GameLogic.scala 258:39]
  reg [10:0] _T_913; // @[GameLogic.scala 263:43]
  wire [10:0] _T_917 = $signed(_T_913) + 11'sh10; // @[GameLogic.scala 263:59]
  reg [10:0] _T_918; // @[GameLogic.scala 264:43]
  wire  _T_919 = ~btnCReg; // @[GameLogic.scala 267:22]
  wire  _T_920 = shotLoad & _T_919; // @[GameLogic.scala 267:19]
  wire [2:0] _T_923 = $signed(shotCntBig) - 3'sh1; // @[GameLogic.scala 270:32]
  wire  _GEN_890 = _T_920 | _GEN_881; // @[GameLogic.scala 267:32]
  wire  _GEN_893 = _T_920 ? 1'h0 : _GEN_883; // @[GameLogic.scala 267:32]
  wire  _GEN_894 = _T_920 | _GEN_882; // @[GameLogic.scala 267:32]
  wire  _GEN_898 = shotPop_3 ? _GEN_890 : _GEN_881; // @[GameLogic.scala 948:28]
  wire  _GEN_900 = shotPop_3 ? _GEN_893 : _GEN_883; // @[GameLogic.scala 948:28]
  wire  _GEN_901 = shotPop_3 ? _GEN_894 : _GEN_882; // @[GameLogic.scala 948:28]
  wire  _T_924 = $signed(shotCntFast) > 3'sh0; // @[GameLogic.scala 951:44]
  wire  _T_925 = io_sw_2 & _T_924; // @[GameLogic.scala 951:29]
  wire  _T_927 = btnCReg & _T_924; // @[GameLogic.scala 239:18]
  wire  _GEN_902 = _T_927 | shotLoad; // @[GameLogic.scala 239:40]
  reg [10:0] _T_928; // @[GameLogic.scala 244:43]
  wire [10:0] _T_932 = $signed(_T_928) + 11'sh10; // @[GameLogic.scala 244:59]
  reg [10:0] _T_933; // @[GameLogic.scala 245:43]
  wire [2:0] _T_938 = $signed(shotCntFast) - 3'sh1; // @[GameLogic.scala 251:34]
  wire  _GEN_905 = _T_920 | _GEN_884; // @[GameLogic.scala 248:32]
  wire  _GEN_908 = _T_920 ? 1'h0 : _GEN_886; // @[GameLogic.scala 248:32]
  wire  _GEN_909 = _T_920 | _GEN_885; // @[GameLogic.scala 248:32]
  wire  _GEN_913 = shotPop_4 ? _GEN_905 : _GEN_884; // @[GameLogic.scala 953:28]
  wire  _GEN_915 = shotPop_4 ? _GEN_908 : _GEN_886; // @[GameLogic.scala 953:28]
  wire  _GEN_916 = shotPop_4 ? _GEN_909 : _GEN_885; // @[GameLogic.scala 953:28]
  wire  _T_939 = $signed(shotCnt) > 10'sh0; // @[GameLogic.scala 218:29]
  wire  _T_940 = btnCReg & _T_939; // @[GameLogic.scala 218:18]
  wire  _GEN_917 = _T_940 | shotLoad; // @[GameLogic.scala 218:36]
  reg [10:0] _T_941; // @[GameLogic.scala 223:43]
  wire [10:0] _T_945 = $signed(_T_941) + 11'sh10; // @[GameLogic.scala 223:59]
  reg [10:0] _T_946; // @[GameLogic.scala 224:43]
  wire [9:0] _T_951 = $signed(shotCnt) - 10'sh1; // @[GameLogic.scala 230:26]
  wire  _GEN_920 = _T_920 | _GEN_872; // @[GameLogic.scala 227:32]
  wire  _GEN_923 = _T_920 ? 1'h0 : _GEN_874; // @[GameLogic.scala 227:32]
  wire  _GEN_924 = _T_920 | _GEN_873; // @[GameLogic.scala 227:32]
  wire [1:0] _GEN_925 = _T_920 ? 2'h1 : 2'h2; // @[GameLogic.scala 227:32]
  reg [10:0] _T_954; // @[GameLogic.scala 223:43]
  wire [10:0] _T_958 = $signed(_T_954) + 11'sh10; // @[GameLogic.scala 223:59]
  reg [10:0] _T_959; // @[GameLogic.scala 224:43]
  wire  _GEN_929 = _T_920 | _GEN_875; // @[GameLogic.scala 227:32]
  wire  _GEN_932 = _T_920 ? 1'h0 : _GEN_877; // @[GameLogic.scala 227:32]
  wire  _GEN_933 = _T_920 | _GEN_876; // @[GameLogic.scala 227:32]
  reg [10:0] _T_967; // @[GameLogic.scala 223:43]
  wire [10:0] _T_971 = $signed(_T_967) + 11'sh10; // @[GameLogic.scala 223:59]
  reg [10:0] _T_972; // @[GameLogic.scala 224:43]
  wire  _GEN_938 = _T_920 | _GEN_878; // @[GameLogic.scala 227:32]
  wire  _GEN_941 = _T_920 ? 1'h0 : _GEN_880; // @[GameLogic.scala 227:32]
  wire  _GEN_942 = _T_920 | _GEN_879; // @[GameLogic.scala 227:32]
  wire  _GEN_947 = shotPop_2 ? _GEN_938 : _GEN_878; // @[GameLogic.scala 962:34]
  wire  _GEN_949 = shotPop_2 ? _GEN_941 : _GEN_880; // @[GameLogic.scala 962:34]
  wire  _GEN_950 = shotPop_2 ? _GEN_942 : _GEN_879; // @[GameLogic.scala 962:34]
  wire [1:0] _GEN_951 = shotPop_2 ? _GEN_925 : 2'h2; // @[GameLogic.scala 962:34]
  wire  _GEN_955 = shotPop_1 ? _GEN_929 : _GEN_875; // @[GameLogic.scala 960:34]
  wire  _GEN_957 = shotPop_1 ? _GEN_932 : _GEN_877; // @[GameLogic.scala 960:34]
  wire  _GEN_958 = shotPop_1 ? _GEN_933 : _GEN_876; // @[GameLogic.scala 960:34]
  wire [1:0] _GEN_959 = shotPop_1 ? _GEN_925 : _GEN_951; // @[GameLogic.scala 960:34]
  wire  _GEN_962 = shotPop_1 ? _GEN_878 : _GEN_947; // @[GameLogic.scala 960:34]
  wire  _GEN_963 = shotPop_1 ? _GEN_880 : _GEN_949; // @[GameLogic.scala 960:34]
  wire  _GEN_964 = shotPop_1 ? _GEN_879 : _GEN_950; // @[GameLogic.scala 960:34]
  wire  _GEN_968 = shotPop_0 ? _GEN_920 : _GEN_872; // @[GameLogic.scala 958:28]
  wire  _GEN_970 = shotPop_0 ? _GEN_923 : _GEN_874; // @[GameLogic.scala 958:28]
  wire  _GEN_971 = shotPop_0 ? _GEN_924 : _GEN_873; // @[GameLogic.scala 958:28]
  wire [1:0] _GEN_972 = shotPop_0 ? _GEN_925 : _GEN_959; // @[GameLogic.scala 958:28]
  wire  _GEN_975 = shotPop_0 ? _GEN_875 : _GEN_955; // @[GameLogic.scala 958:28]
  wire  _GEN_976 = shotPop_0 ? _GEN_877 : _GEN_957; // @[GameLogic.scala 958:28]
  wire  _GEN_977 = shotPop_0 ? _GEN_876 : _GEN_958; // @[GameLogic.scala 958:28]
  wire  _GEN_980 = shotPop_0 ? _GEN_878 : _GEN_962; // @[GameLogic.scala 958:28]
  wire  _GEN_981 = shotPop_0 ? _GEN_880 : _GEN_963; // @[GameLogic.scala 958:28]
  wire  _GEN_982 = shotPop_0 ? _GEN_879 : _GEN_964; // @[GameLogic.scala 958:28]
  wire  _GEN_987 = _T_925 ? _GEN_913 : _GEN_884; // @[GameLogic.scala 951:51]
  wire  _GEN_989 = _T_925 ? _GEN_915 : _GEN_886; // @[GameLogic.scala 951:51]
  wire  _GEN_990 = _T_925 ? _GEN_916 : _GEN_885; // @[GameLogic.scala 951:51]
  wire  _GEN_993 = _T_925 ? _GEN_872 : _GEN_968; // @[GameLogic.scala 951:51]
  wire  _GEN_995 = _T_925 ? _GEN_874 : _GEN_970; // @[GameLogic.scala 951:51]
  wire  _GEN_996 = _T_925 ? _GEN_873 : _GEN_971; // @[GameLogic.scala 951:51]
  wire [1:0] _GEN_997 = _T_925 ? 2'h2 : _GEN_972; // @[GameLogic.scala 951:51]
  wire  _GEN_1000 = _T_925 ? _GEN_875 : _GEN_975; // @[GameLogic.scala 951:51]
  wire  _GEN_1001 = _T_925 ? _GEN_877 : _GEN_976; // @[GameLogic.scala 951:51]
  wire  _GEN_1002 = _T_925 ? _GEN_876 : _GEN_977; // @[GameLogic.scala 951:51]
  wire  _GEN_1005 = _T_925 ? _GEN_878 : _GEN_980; // @[GameLogic.scala 951:51]
  wire  _GEN_1006 = _T_925 ? _GEN_880 : _GEN_981; // @[GameLogic.scala 951:51]
  wire  _GEN_1007 = _T_925 ? _GEN_879 : _GEN_982; // @[GameLogic.scala 951:51]
  wire  _GEN_1012 = _T_910 ? _GEN_898 : _GEN_881; // @[GameLogic.scala 946:44]
  wire  _GEN_1014 = _T_910 ? _GEN_900 : _GEN_883; // @[GameLogic.scala 946:44]
  wire  _GEN_1015 = _T_910 ? _GEN_901 : _GEN_882; // @[GameLogic.scala 946:44]
  wire  _GEN_1018 = _T_910 ? _GEN_884 : _GEN_987; // @[GameLogic.scala 946:44]
  wire  _GEN_1020 = _T_910 ? _GEN_886 : _GEN_989; // @[GameLogic.scala 946:44]
  wire  _GEN_1021 = _T_910 ? _GEN_885 : _GEN_990; // @[GameLogic.scala 946:44]
  wire  _GEN_1024 = _T_910 ? _GEN_872 : _GEN_993; // @[GameLogic.scala 946:44]
  wire  _GEN_1026 = _T_910 ? _GEN_874 : _GEN_995; // @[GameLogic.scala 946:44]
  wire  _GEN_1027 = _T_910 ? _GEN_873 : _GEN_996; // @[GameLogic.scala 946:44]
  wire [1:0] _GEN_1028 = _T_910 ? 2'h2 : _GEN_997; // @[GameLogic.scala 946:44]
  wire  _GEN_1031 = _T_910 ? _GEN_875 : _GEN_1000; // @[GameLogic.scala 946:44]
  wire  _GEN_1032 = _T_910 ? _GEN_877 : _GEN_1001; // @[GameLogic.scala 946:44]
  wire  _GEN_1033 = _T_910 ? _GEN_876 : _GEN_1002; // @[GameLogic.scala 946:44]
  wire  _GEN_1036 = _T_910 ? _GEN_878 : _GEN_1005; // @[GameLogic.scala 946:44]
  wire  _GEN_1037 = _T_910 ? _GEN_880 : _GEN_1006; // @[GameLogic.scala 946:44]
  wire  _GEN_1038 = _T_910 ? _GEN_879 : _GEN_1007; // @[GameLogic.scala 946:44]
  wire  _GEN_1043 = _T_864 ? _GEN_1012 : _GEN_881; // @[GameLogic.scala 945:22]
  wire  _GEN_1045 = _T_864 ? _GEN_1014 : _GEN_883; // @[GameLogic.scala 945:22]
  wire  _GEN_1046 = _T_864 ? _GEN_1015 : _GEN_882; // @[GameLogic.scala 945:22]
  wire  _GEN_1049 = _T_864 ? _GEN_1018 : _GEN_884; // @[GameLogic.scala 945:22]
  wire  _GEN_1051 = _T_864 ? _GEN_1020 : _GEN_886; // @[GameLogic.scala 945:22]
  wire  _GEN_1052 = _T_864 ? _GEN_1021 : _GEN_885; // @[GameLogic.scala 945:22]
  wire  _GEN_1055 = _T_864 ? _GEN_1024 : _GEN_872; // @[GameLogic.scala 945:22]
  wire  _GEN_1057 = _T_864 ? _GEN_1026 : _GEN_874; // @[GameLogic.scala 945:22]
  wire  _GEN_1058 = _T_864 ? _GEN_1027 : _GEN_873; // @[GameLogic.scala 945:22]
  wire [1:0] _GEN_1059 = _T_864 ? _GEN_1028 : 2'h2; // @[GameLogic.scala 945:22]
  wire  _GEN_1062 = _T_864 ? _GEN_1031 : _GEN_875; // @[GameLogic.scala 945:22]
  wire  _GEN_1063 = _T_864 ? _GEN_1032 : _GEN_877; // @[GameLogic.scala 945:22]
  wire  _GEN_1064 = _T_864 ? _GEN_1033 : _GEN_876; // @[GameLogic.scala 945:22]
  wire  _GEN_1067 = _T_864 ? _GEN_1036 : _GEN_878; // @[GameLogic.scala 945:22]
  wire  _GEN_1068 = _T_864 ? _GEN_1037 : _GEN_880; // @[GameLogic.scala 945:22]
  wire  _GEN_1069 = _T_864 ? _GEN_1038 : _GEN_879; // @[GameLogic.scala 945:22]
  wire  _T_978 = 4'hc == stateReg; // @[Conditional.scala 37:30]
  reg  _T_979; // @[GameLogic.scala 128:23]
  reg  _T_980; // @[GameLogic.scala 129:23]
  reg [2:0] _T_981; // @[GameLogic.scala 131:25]
  reg [2:0] _T_982; // @[GameLogic.scala 132:25]
  reg [2:0] _T_983; // @[GameLogic.scala 133:25]
  wire  _T_984 = $signed(Xstart_125) > 11'sh2a0; // @[GameLogic.scala 135:26]
  wire  _T_985 = $signed(Xstart_126) > 11'sh2a0; // @[GameLogic.scala 138:26]
  wire  _T_986 = $signed(Xstart_127) > 11'sh2a0; // @[GameLogic.scala 141:26]
  wire [4:0] _GEN_4462 = {{2{_T_981[2]}},_T_981}; // @[GameLogic.scala 144:35]
  wire [4:0] _T_989 = 5'sha + $signed(_GEN_4462); // @[GameLogic.scala 144:35]
  wire [10:0] _GEN_4463 = {{6{_T_989[4]}},_T_989}; // @[GameLogic.scala 122:44]
  wire [10:0] _T_992 = $signed(Xstart_125) - $signed(_GEN_4463); // @[GameLogic.scala 122:44]
  wire  _T_993 = $signed(Xstart_125) <= 11'sh2; // @[GameLogic.scala 109:28]
  wire  _T_998 = $signed(Randomizer_35_io_out) <= 6'sh8; // @[GameLogic.scala 113:27]
  wire  _T_999 = $signed(Xstart_125) <= 11'sh160; // @[GameLogic.scala 146:26]
  wire  _GEN_1078 = _T_999 | _T_979; // @[GameLogic.scala 146:38]
  wire  _T_1000 = $signed(Xstart_126) <= 11'sh160; // @[GameLogic.scala 149:26]
  wire  _GEN_1079 = _T_1000 | _T_980; // @[GameLogic.scala 149:38]
  wire [4:0] _GEN_4465 = {{2{_T_982[2]}},_T_982}; // @[GameLogic.scala 153:36]
  wire [4:0] _T_1004 = 5'sh8 + $signed(_GEN_4465); // @[GameLogic.scala 153:36]
  wire [10:0] _GEN_4466 = {{6{_T_1004[4]}},_T_1004}; // @[GameLogic.scala 122:44]
  wire [10:0] _T_1007 = $signed(Xstart_126) - $signed(_GEN_4466); // @[GameLogic.scala 122:44]
  wire  _T_1008 = $signed(Xstart_126) <= 11'sh2; // @[GameLogic.scala 109:28]
  wire  _T_1013 = $signed(Randomizer_37_io_out) <= 6'sh8; // @[GameLogic.scala 113:27]
  wire [3:0] _GEN_4468 = {{1{_T_983[2]}},_T_983}; // @[GameLogic.scala 156:36]
  wire [3:0] _T_1017 = 4'sh6 + $signed(_GEN_4468); // @[GameLogic.scala 156:36]
  wire [10:0] _GEN_4469 = {{7{_T_1017[3]}},_T_1017}; // @[GameLogic.scala 122:44]
  wire [10:0] _T_1020 = $signed(Xstart_127) - $signed(_GEN_4469); // @[GameLogic.scala 122:44]
  wire  _T_1021 = $signed(Xstart_127) <= 11'sh2; // @[GameLogic.scala 109:28]
  wire  _T_1026 = $signed(Randomizer_39_io_out) <= 6'sh8; // @[GameLogic.scala 113:27]
  wire  _T_1027 = $signed(cnt) == 10'sh5; // @[GameLogic.scala 973:16]
  wire  _T_1028 = count5 == 8'h1; // @[GameLogic.scala 976:19]
  reg  _T_1029; // @[GameLogic.scala 128:23]
  reg  _T_1030; // @[GameLogic.scala 129:23]
  reg [2:0] _T_1031; // @[GameLogic.scala 131:25]
  reg [2:0] _T_1032; // @[GameLogic.scala 132:25]
  reg [2:0] _T_1033; // @[GameLogic.scala 133:25]
  wire  _T_1034 = $signed(Xstart_122) > 11'sh2a0; // @[GameLogic.scala 135:26]
  wire  _T_1035 = $signed(Xstart_123) > 11'sh2a0; // @[GameLogic.scala 138:26]
  wire  _T_1036 = $signed(Xstart_124) > 11'sh2a0; // @[GameLogic.scala 141:26]
  wire [4:0] _GEN_4471 = {{2{_T_1031[2]}},_T_1031}; // @[GameLogic.scala 144:35]
  wire [4:0] _T_1039 = 5'sha + $signed(_GEN_4471); // @[GameLogic.scala 144:35]
  wire [10:0] _GEN_4472 = {{6{_T_1039[4]}},_T_1039}; // @[GameLogic.scala 122:44]
  wire [10:0] _T_1042 = $signed(Xstart_122) - $signed(_GEN_4472); // @[GameLogic.scala 122:44]
  wire  _T_1043 = $signed(Xstart_122) <= 11'sh2; // @[GameLogic.scala 109:28]
  wire  _T_1048 = $signed(Randomizer_42_io_out) <= 6'sh8; // @[GameLogic.scala 113:27]
  wire  _T_1049 = $signed(Xstart_122) <= 11'sh160; // @[GameLogic.scala 146:26]
  wire  _GEN_1107 = _T_1049 | _T_1029; // @[GameLogic.scala 146:38]
  wire  _T_1050 = $signed(Xstart_123) <= 11'sh160; // @[GameLogic.scala 149:26]
  wire  _GEN_1108 = _T_1050 | _T_1030; // @[GameLogic.scala 149:38]
  wire [4:0] _GEN_4474 = {{2{_T_1032[2]}},_T_1032}; // @[GameLogic.scala 153:36]
  wire [4:0] _T_1054 = 5'sh8 + $signed(_GEN_4474); // @[GameLogic.scala 153:36]
  wire [10:0] _GEN_4475 = {{6{_T_1054[4]}},_T_1054}; // @[GameLogic.scala 122:44]
  wire [10:0] _T_1057 = $signed(Xstart_123) - $signed(_GEN_4475); // @[GameLogic.scala 122:44]
  wire  _T_1058 = $signed(Xstart_123) <= 11'sh2; // @[GameLogic.scala 109:28]
  wire  _T_1063 = $signed(Randomizer_44_io_out) <= 6'sh8; // @[GameLogic.scala 113:27]
  wire [3:0] _GEN_4477 = {{1{_T_1033[2]}},_T_1033}; // @[GameLogic.scala 156:36]
  wire [3:0] _T_1067 = 4'sh6 + $signed(_GEN_4477); // @[GameLogic.scala 156:36]
  wire [10:0] _GEN_4478 = {{7{_T_1067[3]}},_T_1067}; // @[GameLogic.scala 122:44]
  wire [10:0] _T_1070 = $signed(Xstart_124) - $signed(_GEN_4478); // @[GameLogic.scala 122:44]
  wire  _T_1071 = $signed(Xstart_124) <= 11'sh2; // @[GameLogic.scala 109:28]
  wire  _T_1076 = $signed(Randomizer_46_io_out) <= 6'sh8; // @[GameLogic.scala 113:27]
  wire  _T_1077 = io_btnC | io_btnL; // @[GameLogic.scala 980:28]
  wire  _T_1078 = _T_1077 | io_btnD; // @[GameLogic.scala 980:39]
  wire  _T_1079 = _T_1078 | io_btnU; // @[GameLogic.scala 980:50]
  wire  _T_1080 = _T_1079 | io_btnR; // @[GameLogic.scala 980:61]
  wire  _T_1081 = _T_1080 | start; // @[GameLogic.scala 980:19]
  wire  _T_1083 = $signed(secCnt) <= 8'sh9; // @[GameLogic.scala 981:36]
  wire  _T_1084 = _T_514 & _T_1083; // @[GameLogic.scala 981:26]
  wire  _T_1085 = level == 3'h4; // @[GameLogic.scala 981:52]
  wire  _T_1086 = _T_1084 & _T_1085; // @[GameLogic.scala 981:43]
  wire  _T_1088 = $signed(cnt) == 10'sh3c; // @[GameLogic.scala 992:16]
  wire  _T_1089 = _T_1088 & start; // @[GameLogic.scala 992:25]
  wire [7:0] _T_1092 = $signed(secCnt) + 8'sh1; // @[GameLogic.scala 993:26]
  wire  _T_1093 = $signed(secCnt) == 8'shf; // @[GameLogic.scala 994:35]
  wire  _T_1094 = io_sw_7 & _T_1093; // @[GameLogic.scala 994:25]
  wire  _T_1095 = $signed(secCnt) == 8'sh3c; // @[GameLogic.scala 994:55]
  wire  _T_1096 = _T_1094 | _T_1095; // @[GameLogic.scala 994:45]
  wire  _T_1098 = _T_1096 & _T_864; // @[GameLogic.scala 994:65]
  wire  _T_1100 = _T_1098 & _T_507; // @[GameLogic.scala 994:77]
  wire [2:0] _T_1102 = level + 3'h1; // @[GameLogic.scala 996:26]
  wire  _T_1105 = _T_1095 & _T_1085; // @[GameLogic.scala 999:36]
  wire [3:0] _GEN_1161 = _T_1100 ? 4'h3 : hp; // @[GameLogic.scala 994:93]
  wire  _GEN_1167 = _T_1100 | levelCng; // @[GameLogic.scala 994:93]
  wire [3:0] _GEN_1169 = _T_1089 ? _GEN_1161 : hp; // @[GameLogic.scala 992:35]
  wire [9:0] _T_1109 = $signed(cnt) + 10'sh1; // @[GameLogic.scala 1004:41]
  wire  _T_1112 = cng ? _T_27 : show; // @[GameLogic.scala 1005:18]
  wire  _T_1113 = $signed(cnt) < 10'sh7; // @[GameLogic.scala 1006:21]
  wire  _T_1114 = $signed(cnt) > 10'sh1e; // @[GameLogic.scala 1006:35]
  wire  _T_1115 = $signed(cnt) < 10'sh25; // @[GameLogic.scala 1006:49]
  wire  _T_1116 = _T_1114 & _T_1115; // @[GameLogic.scala 1006:42]
  wire  _T_1117 = _T_1113 | _T_1116; // @[GameLogic.scala 1006:27]
  wire  _T_1119 = cng & _T_282; // @[GameLogic.scala 1007:16]
  wire [3:0] _T_1121 = cngCnt + 4'h1; // @[GameLogic.scala 1008:26]
  wire  _T_1122 = cngCnt >= 4'h5; // @[GameLogic.scala 1009:21]
  wire  _T_1123 = astInteract_0 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1124 = _T_1123 & boxDetection_io_overlap_0_7; // @[GameLogic.scala 1015:50]
  wire  _T_1125 = astInteract_0 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1126 = _T_1125 & boxDetection_io_overlap_2_7; // @[GameLogic.scala 1017:59]
  wire  _T_1127 = astInteract_0 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1128 = _T_1127 & boxDetection_io_overlap_3_7; // @[GameLogic.scala 1017:59]
  wire  _T_1129 = astInteract_0 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1130 = _T_1129 & boxDetection_io_overlap_4_7; // @[GameLogic.scala 1017:59]
  wire  _T_1131 = astInteract_0 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1132 = _T_1131 & boxDetection_io_overlap_5_7; // @[GameLogic.scala 1017:59]
  wire  _T_1133 = astInteract_0 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1134 = _T_1133 & boxDetection_io_overlap_6_7; // @[GameLogic.scala 1017:59]
  wire  _T_1135 = hp > 4'h1; // @[GameLogic.scala 292:15]
  wire [10:0] _GEN_1177 = _T_1135 ? $signed(11'sh40) : $signed(Xstart_0); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1178 = _T_1135 ? $signed(11'she0) : $signed(Ystart_0); // @[GameLogic.scala 292:22]
  wire  _T_1137 = shipInteract & _T_864; // @[GameLogic.scala 297:25]
  wire [3:0] _T_1139 = hp - 4'h1; // @[GameLogic.scala 298:18]
  wire [3:0] _GEN_1179 = _T_1137 ? _T_1139 : _GEN_1169; // @[GameLogic.scala 297:38]
  wire  _GEN_1181 = _T_1137 ? 1'h0 : shipInteract; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1182 = die_0 ? $signed(_GEN_1177) : $signed(Xstart_0); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1183 = die_0 ? $signed(_GEN_1178) : $signed(Ystart_0); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1184 = die_0 ? _GEN_1179 : _GEN_1169; // @[GameLogic.scala 286:18]
  wire  _GEN_1186 = die_0 ? _GEN_1181 : shipInteract; // @[GameLogic.scala 286:18]
  wire  _T_1140 = astInteract_1 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1141 = _T_1140 & boxDetection_io_overlap_0_8; // @[GameLogic.scala 1015:50]
  wire  _T_1142 = astInteract_1 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1143 = _T_1142 & boxDetection_io_overlap_2_8; // @[GameLogic.scala 1017:59]
  wire  _T_1144 = astInteract_1 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1145 = _T_1144 & boxDetection_io_overlap_3_8; // @[GameLogic.scala 1017:59]
  wire  _T_1146 = astInteract_1 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1147 = _T_1146 & boxDetection_io_overlap_4_8; // @[GameLogic.scala 1017:59]
  wire  _T_1148 = astInteract_1 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1149 = _T_1148 & boxDetection_io_overlap_5_8; // @[GameLogic.scala 1017:59]
  wire  _T_1150 = astInteract_1 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1151 = _T_1150 & boxDetection_io_overlap_6_8; // @[GameLogic.scala 1017:59]
  wire [10:0] _GEN_1187 = _T_1135 ? $signed(11'sh40) : $signed(_GEN_1182); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1188 = _T_1135 ? $signed(11'she0) : $signed(_GEN_1183); // @[GameLogic.scala 292:22]
  wire [3:0] _GEN_1189 = _T_1137 ? _T_1139 : _GEN_1184; // @[GameLogic.scala 297:38]
  wire  _GEN_1191 = _T_1137 ? 1'h0 : _GEN_1186; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1192 = die_1 ? $signed(_GEN_1187) : $signed(_GEN_1182); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1193 = die_1 ? $signed(_GEN_1188) : $signed(_GEN_1183); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1194 = die_1 ? _GEN_1189 : _GEN_1184; // @[GameLogic.scala 286:18]
  wire  _GEN_1196 = die_1 ? _GEN_1191 : _GEN_1186; // @[GameLogic.scala 286:18]
  wire  _T_1157 = astInteract_2 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1158 = _T_1157 & boxDetection_io_overlap_0_9; // @[GameLogic.scala 1015:50]
  wire  _T_1159 = astInteract_2 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1160 = _T_1159 & boxDetection_io_overlap_2_9; // @[GameLogic.scala 1017:59]
  wire  _T_1161 = astInteract_2 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1162 = _T_1161 & boxDetection_io_overlap_3_9; // @[GameLogic.scala 1017:59]
  wire  _T_1163 = astInteract_2 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1164 = _T_1163 & boxDetection_io_overlap_4_9; // @[GameLogic.scala 1017:59]
  wire  _T_1165 = astInteract_2 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1166 = _T_1165 & boxDetection_io_overlap_5_9; // @[GameLogic.scala 1017:59]
  wire  _T_1167 = astInteract_2 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1168 = _T_1167 & boxDetection_io_overlap_6_9; // @[GameLogic.scala 1017:59]
  wire [10:0] _GEN_1197 = _T_1135 ? $signed(11'sh40) : $signed(_GEN_1192); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1198 = _T_1135 ? $signed(11'she0) : $signed(_GEN_1193); // @[GameLogic.scala 292:22]
  wire [3:0] _GEN_1199 = _T_1137 ? _T_1139 : _GEN_1194; // @[GameLogic.scala 297:38]
  wire  _GEN_1201 = _T_1137 ? 1'h0 : _GEN_1196; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1202 = die_2 ? $signed(_GEN_1197) : $signed(_GEN_1192); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1203 = die_2 ? $signed(_GEN_1198) : $signed(_GEN_1193); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1204 = die_2 ? _GEN_1199 : _GEN_1194; // @[GameLogic.scala 286:18]
  wire  _GEN_1206 = die_2 ? _GEN_1201 : _GEN_1196; // @[GameLogic.scala 286:18]
  wire  _T_1174 = astInteract_3 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1175 = _T_1174 & boxDetection_io_overlap_0_10; // @[GameLogic.scala 1015:50]
  wire  _T_1176 = astInteract_3 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1177 = _T_1176 & boxDetection_io_overlap_2_10; // @[GameLogic.scala 1017:59]
  wire  _T_1178 = astInteract_3 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1179 = _T_1178 & boxDetection_io_overlap_3_10; // @[GameLogic.scala 1017:59]
  wire  _T_1180 = astInteract_3 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1181 = _T_1180 & boxDetection_io_overlap_4_10; // @[GameLogic.scala 1017:59]
  wire  _T_1182 = astInteract_3 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1183 = _T_1182 & boxDetection_io_overlap_5_10; // @[GameLogic.scala 1017:59]
  wire  _T_1184 = astInteract_3 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1185 = _T_1184 & boxDetection_io_overlap_6_10; // @[GameLogic.scala 1017:59]
  wire [10:0] _GEN_1207 = _T_1135 ? $signed(11'sh40) : $signed(_GEN_1202); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1208 = _T_1135 ? $signed(11'she0) : $signed(_GEN_1203); // @[GameLogic.scala 292:22]
  wire [3:0] _GEN_1209 = _T_1137 ? _T_1139 : _GEN_1204; // @[GameLogic.scala 297:38]
  wire  _GEN_1211 = _T_1137 ? 1'h0 : _GEN_1206; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1212 = die_3 ? $signed(_GEN_1207) : $signed(_GEN_1202); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1213 = die_3 ? $signed(_GEN_1208) : $signed(_GEN_1203); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1214 = die_3 ? _GEN_1209 : _GEN_1204; // @[GameLogic.scala 286:18]
  wire  _GEN_1216 = die_3 ? _GEN_1211 : _GEN_1206; // @[GameLogic.scala 286:18]
  wire  _T_1191 = astInteract_4 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1192 = _T_1191 & boxDetection_io_overlap_0_11; // @[GameLogic.scala 1015:50]
  wire  _T_1193 = astInteract_4 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1194 = _T_1193 & boxDetection_io_overlap_2_11; // @[GameLogic.scala 1017:59]
  wire  _T_1195 = astInteract_4 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1196 = _T_1195 & boxDetection_io_overlap_3_11; // @[GameLogic.scala 1017:59]
  wire  _T_1197 = astInteract_4 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1198 = _T_1197 & boxDetection_io_overlap_4_11; // @[GameLogic.scala 1017:59]
  wire  _T_1199 = astInteract_4 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1200 = _T_1199 & boxDetection_io_overlap_5_11; // @[GameLogic.scala 1017:59]
  wire  _T_1201 = astInteract_4 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1202 = _T_1201 & boxDetection_io_overlap_6_11; // @[GameLogic.scala 1017:59]
  wire [10:0] _GEN_1217 = _T_1135 ? $signed(11'sh40) : $signed(_GEN_1212); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1218 = _T_1135 ? $signed(11'she0) : $signed(_GEN_1213); // @[GameLogic.scala 292:22]
  wire [3:0] _GEN_1219 = _T_1137 ? _T_1139 : _GEN_1214; // @[GameLogic.scala 297:38]
  wire  _GEN_1221 = _T_1137 ? 1'h0 : _GEN_1216; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1222 = die_4 ? $signed(_GEN_1217) : $signed(_GEN_1212); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1223 = die_4 ? $signed(_GEN_1218) : $signed(_GEN_1213); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1224 = die_4 ? _GEN_1219 : _GEN_1214; // @[GameLogic.scala 286:18]
  wire  _GEN_1226 = die_4 ? _GEN_1221 : _GEN_1216; // @[GameLogic.scala 286:18]
  wire  _T_1208 = astInteract_5 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1209 = _T_1208 & boxDetection_io_overlap_0_12; // @[GameLogic.scala 1015:50]
  wire  _T_1210 = astInteract_5 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1211 = _T_1210 & boxDetection_io_overlap_2_12; // @[GameLogic.scala 1017:59]
  wire  _T_1212 = astInteract_5 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1213 = _T_1212 & boxDetection_io_overlap_3_12; // @[GameLogic.scala 1017:59]
  wire  _T_1214 = astInteract_5 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1215 = _T_1214 & boxDetection_io_overlap_4_12; // @[GameLogic.scala 1017:59]
  wire  _T_1216 = astInteract_5 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1217 = _T_1216 & boxDetection_io_overlap_5_12; // @[GameLogic.scala 1017:59]
  wire  _T_1218 = astInteract_5 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1219 = _T_1218 & boxDetection_io_overlap_6_12; // @[GameLogic.scala 1017:59]
  wire [10:0] _GEN_1227 = _T_1135 ? $signed(11'sh40) : $signed(_GEN_1222); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1228 = _T_1135 ? $signed(11'she0) : $signed(_GEN_1223); // @[GameLogic.scala 292:22]
  wire [3:0] _GEN_1229 = _T_1137 ? _T_1139 : _GEN_1224; // @[GameLogic.scala 297:38]
  wire  _GEN_1231 = _T_1137 ? 1'h0 : _GEN_1226; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1232 = die_5 ? $signed(_GEN_1227) : $signed(_GEN_1222); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1233 = die_5 ? $signed(_GEN_1228) : $signed(_GEN_1223); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1234 = die_5 ? _GEN_1229 : _GEN_1224; // @[GameLogic.scala 286:18]
  wire  _GEN_1236 = die_5 ? _GEN_1231 : _GEN_1226; // @[GameLogic.scala 286:18]
  wire  _T_1225 = astInteract_6 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1226 = _T_1225 & boxDetection_io_overlap_0_13; // @[GameLogic.scala 1015:50]
  wire  _T_1227 = astInteract_6 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1228 = _T_1227 & boxDetection_io_overlap_2_13; // @[GameLogic.scala 1017:59]
  wire  _T_1229 = astInteract_6 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1230 = _T_1229 & boxDetection_io_overlap_3_13; // @[GameLogic.scala 1017:59]
  wire  _T_1231 = astInteract_6 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1232 = _T_1231 & boxDetection_io_overlap_4_13; // @[GameLogic.scala 1017:59]
  wire  _T_1233 = astInteract_6 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1234 = _T_1233 & boxDetection_io_overlap_5_13; // @[GameLogic.scala 1017:59]
  wire  _T_1235 = astInteract_6 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1236 = _T_1235 & boxDetection_io_overlap_6_13; // @[GameLogic.scala 1017:59]
  wire [10:0] _GEN_1237 = _T_1135 ? $signed(11'sh40) : $signed(_GEN_1232); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1238 = _T_1135 ? $signed(11'she0) : $signed(_GEN_1233); // @[GameLogic.scala 292:22]
  wire [3:0] _GEN_1239 = _T_1137 ? _T_1139 : _GEN_1234; // @[GameLogic.scala 297:38]
  wire  _GEN_1241 = _T_1137 ? 1'h0 : _GEN_1236; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1242 = die_6 ? $signed(_GEN_1237) : $signed(_GEN_1232); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1243 = die_6 ? $signed(_GEN_1238) : $signed(_GEN_1233); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1244 = die_6 ? _GEN_1239 : _GEN_1234; // @[GameLogic.scala 286:18]
  wire  _GEN_1246 = die_6 ? _GEN_1241 : _GEN_1236; // @[GameLogic.scala 286:18]
  wire  _T_1242 = astInteract_7 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1243 = _T_1242 & boxDetection_io_overlap_0_14; // @[GameLogic.scala 1015:50]
  wire  _T_1244 = astInteract_7 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1245 = _T_1244 & boxDetection_io_overlap_2_14; // @[GameLogic.scala 1017:59]
  wire  _T_1246 = astInteract_7 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1247 = _T_1246 & boxDetection_io_overlap_3_14; // @[GameLogic.scala 1017:59]
  wire  _T_1248 = astInteract_7 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1249 = _T_1248 & boxDetection_io_overlap_4_14; // @[GameLogic.scala 1017:59]
  wire  _T_1250 = astInteract_7 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1251 = _T_1250 & boxDetection_io_overlap_5_14; // @[GameLogic.scala 1017:59]
  wire  _T_1252 = astInteract_7 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1253 = _T_1252 & boxDetection_io_overlap_6_14; // @[GameLogic.scala 1017:59]
  wire [10:0] _GEN_1247 = _T_1135 ? $signed(11'sh40) : $signed(_GEN_1242); // @[GameLogic.scala 292:22]
  wire [10:0] _GEN_1248 = _T_1135 ? $signed(11'she0) : $signed(_GEN_1243); // @[GameLogic.scala 292:22]
  wire [3:0] _GEN_1249 = _T_1137 ? _T_1139 : _GEN_1244; // @[GameLogic.scala 297:38]
  wire  _GEN_1251 = _T_1137 ? 1'h0 : _GEN_1246; // @[GameLogic.scala 297:38]
  wire [10:0] _GEN_1252 = die_7 ? $signed(_GEN_1247) : $signed(_GEN_1242); // @[GameLogic.scala 286:18]
  wire [10:0] _GEN_1253 = die_7 ? $signed(_GEN_1248) : $signed(_GEN_1243); // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1254 = die_7 ? _GEN_1249 : _GEN_1244; // @[GameLogic.scala 286:18]
  wire  _GEN_1256 = die_7 ? _GEN_1251 : _GEN_1246; // @[GameLogic.scala 286:18]
  wire  _T_1259 = astInteract_8 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1260 = _T_1259 & boxDetection_io_overlap_0_15; // @[GameLogic.scala 1015:50]
  wire  _T_1261 = astInteract_8 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1262 = _T_1261 & boxDetection_io_overlap_2_15; // @[GameLogic.scala 1017:59]
  wire  _T_1263 = astInteract_8 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1264 = _T_1263 & boxDetection_io_overlap_3_15; // @[GameLogic.scala 1017:59]
  wire  _T_1265 = astInteract_8 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1266 = _T_1265 & boxDetection_io_overlap_4_15; // @[GameLogic.scala 1017:59]
  wire  _T_1267 = astInteract_8 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1268 = _T_1267 & boxDetection_io_overlap_5_15; // @[GameLogic.scala 1017:59]
  wire  _T_1269 = astInteract_8 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1270 = _T_1269 & boxDetection_io_overlap_6_15; // @[GameLogic.scala 1017:59]
  wire  _GEN_1261 = _T_1137 ? 1'h0 : _GEN_1256; // @[GameLogic.scala 297:38]
  wire  _GEN_1266 = die_8 ? _GEN_1261 : _GEN_1256; // @[GameLogic.scala 286:18]
  wire  _T_1276 = astInteract_9 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1277 = _T_1276 & boxDetection_io_overlap_0_16; // @[GameLogic.scala 1015:50]
  wire  _T_1278 = astInteract_9 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1279 = _T_1278 & boxDetection_io_overlap_2_16; // @[GameLogic.scala 1017:59]
  wire  _T_1280 = astInteract_9 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1281 = _T_1280 & boxDetection_io_overlap_3_16; // @[GameLogic.scala 1017:59]
  wire  _T_1282 = astInteract_9 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1283 = _T_1282 & boxDetection_io_overlap_4_16; // @[GameLogic.scala 1017:59]
  wire  _T_1284 = astInteract_9 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1285 = _T_1284 & boxDetection_io_overlap_5_16; // @[GameLogic.scala 1017:59]
  wire  _GEN_1271 = _T_1137 ? 1'h0 : _GEN_1266; // @[GameLogic.scala 297:38]
  wire  _GEN_1276 = die_9 ? _GEN_1271 : _GEN_1266; // @[GameLogic.scala 286:18]
  wire  _T_1293 = astInteract_10 & shipInteract; // @[GameLogic.scala 1015:34]
  wire  _T_1294 = _T_1293 & boxDetection_io_overlap_0_17; // @[GameLogic.scala 1015:50]
  wire  _T_1295 = astInteract_10 & shotInteract_0; // @[GameLogic.scala 1017:40]
  wire  _T_1296 = _T_1295 & boxDetection_io_overlap_2_17; // @[GameLogic.scala 1017:59]
  wire  _T_1297 = astInteract_10 & shotInteract_1; // @[GameLogic.scala 1017:40]
  wire  _T_1298 = _T_1297 & boxDetection_io_overlap_3_17; // @[GameLogic.scala 1017:59]
  wire  _T_1299 = astInteract_10 & shotInteract_2; // @[GameLogic.scala 1017:40]
  wire  _T_1300 = _T_1299 & boxDetection_io_overlap_4_17; // @[GameLogic.scala 1017:59]
  wire  _T_1301 = astInteract_10 & shotInteract_3; // @[GameLogic.scala 1017:40]
  wire  _T_1302 = _T_1301 & boxDetection_io_overlap_5_17; // @[GameLogic.scala 1017:59]
  wire  _T_1303 = astInteract_10 & shotInteract_4; // @[GameLogic.scala 1017:40]
  wire  _T_1304 = _T_1303 & boxDetection_io_overlap_6_17; // @[GameLogic.scala 1017:59]
  wire  _GEN_1281 = _T_1137 ? 1'h0 : _GEN_1276; // @[GameLogic.scala 297:38]
  wire  _GEN_1286 = die_10 ? _GEN_1281 : _GEN_1276; // @[GameLogic.scala 286:18]
  wire  _T_1311 = cng & _T_28; // @[GameLogic.scala 1021:16]
  wire [5:0] _T_1314 = $signed(spwnProt) + 6'sh1; // @[GameLogic.scala 1022:30]
  wire  _T_1315 = $signed(spwnProt) >= 6'sh6; // @[GameLogic.scala 1024:21]
  wire  _GEN_1288 = _T_1315 | _GEN_1286; // @[GameLogic.scala 1024:29]
  wire  _GEN_1294 = io_sw_0 | _T_1081; // @[GameLogic.scala 1028:22]
  wire  _T_1360 = $signed(shotCntFast) > 3'sh1; // @[GameLogic.scala 327:47]
  wire  _T_1361 = $signed(shotCntBig) > 3'sh1; // @[GameLogic.scala 328:46]
  wire  _T_1362 = $signed(shotCnt) > 10'sh5; // @[GameLogic.scala 329:43]
  wire  _T_1364 = $signed(shotCntFast) > 3'sh2; // @[GameLogic.scala 327:47]
  wire  _T_1365 = $signed(shotCntBig) > 3'sh2; // @[GameLogic.scala 328:46]
  wire  _T_1366 = $signed(shotCnt) > 10'sha; // @[GameLogic.scala 329:43]
  wire  _T_1367 = hp > 4'h2; // @[GameLogic.scala 330:38]
  wire [5:0] _T_1368 = 5'sh8 * 5'sh0; // @[GameLogic.scala 335:55]
  wire [6:0] _T_1369 = {{1{_T_1368[5]}},_T_1368}; // @[GameLogic.scala 335:48]
  wire [5:0] _T_1371 = _T_1369[5:0]; // @[GameLogic.scala 335:48]
  wire [7:0] _GEN_4480 = {{2{_T_1371[5]}},_T_1371}; // @[GameLogic.scala 335:42]
  wire  _T_1372 = $signed(secCnt) > $signed(_GEN_4480); // @[GameLogic.scala 335:42]
  wire [5:0] _T_1376 = 6'sh8 + $signed(_T_1368); // @[GameLogic.scala 335:79]
  wire [7:0] _GEN_4481 = {{2{_T_1376[5]}},_T_1376}; // @[GameLogic.scala 335:72]
  wire  _T_1377 = $signed(secCnt) <= $signed(_GEN_4481); // @[GameLogic.scala 335:72]
  wire  _T_1378 = _T_1372 & _T_1377; // @[GameLogic.scala 335:62]
  wire [6:0] _T_1379 = 5'sh8 * 5'sh1; // @[GameLogic.scala 335:55]
  wire [7:0] _T_1380 = {{1{_T_1379[6]}},_T_1379}; // @[GameLogic.scala 335:48]
  wire [6:0] _T_1382 = _T_1380[6:0]; // @[GameLogic.scala 335:48]
  wire [7:0] _GEN_4482 = {{1{_T_1382[6]}},_T_1382}; // @[GameLogic.scala 335:42]
  wire  _T_1383 = $signed(secCnt) > $signed(_GEN_4482); // @[GameLogic.scala 335:42]
  wire [6:0] _T_1387 = 7'sh8 + $signed(_T_1379); // @[GameLogic.scala 335:79]
  wire [7:0] _GEN_4483 = {{1{_T_1387[6]}},_T_1387}; // @[GameLogic.scala 335:72]
  wire  _T_1388 = $signed(secCnt) <= $signed(_GEN_4483); // @[GameLogic.scala 335:72]
  wire  _T_1389 = _T_1383 & _T_1388; // @[GameLogic.scala 335:62]
  wire [7:0] _T_1390 = 5'sh8 * 5'sh2; // @[GameLogic.scala 335:55]
  wire [8:0] _T_1391 = {{1{_T_1390[7]}},_T_1390}; // @[GameLogic.scala 335:48]
  wire [7:0] _T_1393 = _T_1391[7:0]; // @[GameLogic.scala 335:48]
  wire  _T_1394 = $signed(secCnt) > $signed(_T_1393); // @[GameLogic.scala 335:42]
  wire [7:0] _T_1398 = 8'sh8 + $signed(_T_1390); // @[GameLogic.scala 335:79]
  wire  _T_1399 = $signed(secCnt) <= $signed(_T_1398); // @[GameLogic.scala 335:72]
  wire  _T_1400 = _T_1394 & _T_1399; // @[GameLogic.scala 335:62]
  wire [7:0] _T_1401 = 5'sh8 * 5'sh3; // @[GameLogic.scala 335:55]
  wire [8:0] _T_1402 = {{1{_T_1401[7]}},_T_1401}; // @[GameLogic.scala 335:48]
  wire [7:0] _T_1404 = _T_1402[7:0]; // @[GameLogic.scala 335:48]
  wire  _T_1405 = $signed(secCnt) > $signed(_T_1404); // @[GameLogic.scala 335:42]
  wire [7:0] _T_1409 = 8'sh8 + $signed(_T_1401); // @[GameLogic.scala 335:79]
  wire  _T_1410 = $signed(secCnt) <= $signed(_T_1409); // @[GameLogic.scala 335:72]
  wire  _T_1411 = _T_1405 & _T_1410; // @[GameLogic.scala 335:62]
  wire [8:0] _T_1412 = 5'sh8 * 5'sh4; // @[GameLogic.scala 335:55]
  wire [9:0] _T_1413 = {{1{_T_1412[8]}},_T_1412}; // @[GameLogic.scala 335:48]
  wire [8:0] _T_1415 = _T_1413[8:0]; // @[GameLogic.scala 335:48]
  wire [8:0] _GEN_4484 = {{1{secCnt[7]}},secCnt}; // @[GameLogic.scala 335:42]
  wire  _T_1416 = $signed(_GEN_4484) > $signed(_T_1415); // @[GameLogic.scala 335:42]
  wire [8:0] _T_1420 = 9'sh8 + $signed(_T_1412); // @[GameLogic.scala 335:79]
  wire  _T_1421 = $signed(_GEN_4484) <= $signed(_T_1420); // @[GameLogic.scala 335:72]
  wire  _T_1422 = _T_1416 & _T_1421; // @[GameLogic.scala 335:62]
  wire [8:0] _T_1423 = 5'sh8 * 5'sh5; // @[GameLogic.scala 335:55]
  wire [9:0] _T_1424 = {{1{_T_1423[8]}},_T_1423}; // @[GameLogic.scala 335:48]
  wire [8:0] _T_1426 = _T_1424[8:0]; // @[GameLogic.scala 335:48]
  wire  _T_1427 = $signed(_GEN_4484) > $signed(_T_1426); // @[GameLogic.scala 335:42]
  wire [8:0] _T_1431 = 9'sh8 + $signed(_T_1423); // @[GameLogic.scala 335:79]
  wire  _T_1432 = $signed(_GEN_4484) <= $signed(_T_1431); // @[GameLogic.scala 335:72]
  wire  _T_1433 = _T_1427 & _T_1432; // @[GameLogic.scala 335:62]
  wire [8:0] _T_1434 = 5'sh8 * 5'sh6; // @[GameLogic.scala 335:55]
  wire [9:0] _T_1435 = {{1{_T_1434[8]}},_T_1434}; // @[GameLogic.scala 335:48]
  wire [8:0] _T_1437 = _T_1435[8:0]; // @[GameLogic.scala 335:48]
  wire  _T_1438 = $signed(_GEN_4484) > $signed(_T_1437); // @[GameLogic.scala 335:42]
  wire [8:0] _T_1442 = 9'sh8 + $signed(_T_1434); // @[GameLogic.scala 335:79]
  wire  _T_1443 = $signed(_GEN_4484) <= $signed(_T_1442); // @[GameLogic.scala 335:72]
  wire  _T_1444 = _T_1438 & _T_1443; // @[GameLogic.scala 335:62]
  wire [8:0] _T_1445 = 5'sh8 * 5'sh7; // @[GameLogic.scala 335:55]
  wire [9:0] _T_1446 = {{1{_T_1445[8]}},_T_1445}; // @[GameLogic.scala 335:48]
  wire [8:0] _T_1448 = _T_1446[8:0]; // @[GameLogic.scala 335:48]
  wire  _T_1449 = $signed(_GEN_4484) > $signed(_T_1448); // @[GameLogic.scala 335:42]
  wire [8:0] _T_1453 = 9'sh8 + $signed(_T_1445); // @[GameLogic.scala 335:79]
  wire  _T_1454 = $signed(_GEN_4484) <= $signed(_T_1453); // @[GameLogic.scala 335:72]
  wire  _T_1455 = _T_1449 & _T_1454; // @[GameLogic.scala 335:62]
  wire  _T_1456 = 4'hd == stateReg; // @[Conditional.scala 37:30]
  wire  _GEN_1352 = _T_978 ? _T_1112 : show; // @[Conditional.scala 39:67]
  wire  _GEN_1363 = _T_978 ? _GEN_1288 : shipInteract; // @[Conditional.scala 39:67]
  wire  _GEN_1427 = _T_978 ? _T_282 : spriteVisibleReg_26; // @[Conditional.scala 39:67]
  wire  _GEN_1430 = _T_978 ? _T_501 : spriteVisibleReg_30; // @[Conditional.scala 39:67]
  wire  _GEN_1433 = _T_978 ? _T_282 : spriteVisibleReg_27; // @[Conditional.scala 39:67]
  wire  _GEN_1436 = _T_978 ? _T_501 : spriteVisibleReg_31; // @[Conditional.scala 39:67]
  wire  _GEN_1439 = _T_978 ? _T_282 : spriteVisibleReg_28; // @[Conditional.scala 39:67]
  wire  _GEN_1442 = _T_978 ? _T_501 : spriteVisibleReg_32; // @[Conditional.scala 39:67]
  wire  _GEN_1445 = _T_978 ? _T_282 : spriteVisibleReg_29; // @[Conditional.scala 39:67]
  wire  _GEN_1448 = _T_978 ? _T_501 : spriteVisibleReg_33; // @[Conditional.scala 39:67]
  wire  _GEN_1451 = _T_978 ? _T_924 : spriteVisibleReg_72; // @[Conditional.scala 39:67]
  wire  _GEN_1452 = _T_978 ? _T_909 : spriteVisibleReg_66; // @[Conditional.scala 39:67]
  wire  _GEN_1453 = _T_978 ? _T_939 : spriteVisibleReg_57; // @[Conditional.scala 39:67]
  wire  _GEN_1454 = _T_978 ? _T_864 : spriteVisibleReg_61; // @[Conditional.scala 39:67]
  wire  _GEN_1455 = _T_978 ? _T_1360 : spriteVisibleReg_71; // @[Conditional.scala 39:67]
  wire  _GEN_1456 = _T_978 ? _T_1361 : spriteVisibleReg_65; // @[Conditional.scala 39:67]
  wire  _GEN_1457 = _T_978 ? _T_1362 : spriteVisibleReg_56; // @[Conditional.scala 39:67]
  wire  _GEN_1458 = _T_978 ? _T_1135 : spriteVisibleReg_62; // @[Conditional.scala 39:67]
  wire  _GEN_1459 = _T_978 ? _T_1364 : spriteVisibleReg_70; // @[Conditional.scala 39:67]
  wire  _GEN_1460 = _T_978 ? _T_1365 : spriteVisibleReg_64; // @[Conditional.scala 39:67]
  wire  _GEN_1461 = _T_978 ? _T_1366 : spriteVisibleReg_55; // @[Conditional.scala 39:67]
  wire  _GEN_1462 = _T_978 ? _T_1367 : spriteVisibleReg_63; // @[Conditional.scala 39:67]
  wire  _GEN_1463 = _T_978 ? _T_1378 : spriteVisibleReg_44; // @[Conditional.scala 39:67]
  wire  _GEN_1466 = _T_978 ? _T_1389 : spriteVisibleReg_45; // @[Conditional.scala 39:67]
  wire  _GEN_1469 = _T_978 ? _T_1400 : spriteVisibleReg_46; // @[Conditional.scala 39:67]
  wire  _GEN_1472 = _T_978 ? _T_1411 : spriteVisibleReg_47; // @[Conditional.scala 39:67]
  wire  _GEN_1475 = _T_978 ? _T_1422 : spriteVisibleReg_48; // @[Conditional.scala 39:67]
  wire  _GEN_1478 = _T_978 ? _T_1433 : spriteVisibleReg_49; // @[Conditional.scala 39:67]
  wire  _GEN_1481 = _T_978 ? _T_1444 : spriteVisibleReg_50; // @[Conditional.scala 39:67]
  wire  _GEN_1484 = _T_978 ? _T_1455 : spriteVisibleReg_51; // @[Conditional.scala 39:67]
  wire  _GEN_1488 = _T_978 ? 1'h0 : _T_1456; // @[Conditional.scala 39:67]
  wire  _GEN_1490 = _T_887 ? _GEN_1055 : spriteVisibleReg_2; // @[Conditional.scala 39:67]
  wire  _GEN_1491 = _T_887 ? _GEN_1058 : shotInteract_0; // @[Conditional.scala 39:67]
  wire  _GEN_1492 = _T_887 ? _GEN_1057 : shotPop_0; // @[Conditional.scala 39:67]
  wire  _GEN_1494 = _T_887 ? _GEN_1062 : spriteVisibleReg_3; // @[Conditional.scala 39:67]
  wire  _GEN_1495 = _T_887 ? _GEN_1064 : shotInteract_1; // @[Conditional.scala 39:67]
  wire  _GEN_1496 = _T_887 ? _GEN_1063 : shotPop_1; // @[Conditional.scala 39:67]
  wire  _GEN_1498 = _T_887 ? _GEN_1067 : spriteVisibleReg_4; // @[Conditional.scala 39:67]
  wire  _GEN_1499 = _T_887 ? _GEN_1069 : shotInteract_2; // @[Conditional.scala 39:67]
  wire  _GEN_1500 = _T_887 ? _GEN_1068 : shotPop_2; // @[Conditional.scala 39:67]
  wire  _GEN_1502 = _T_887 ? _GEN_1043 : spriteVisibleReg_5; // @[Conditional.scala 39:67]
  wire  _GEN_1503 = _T_887 ? _GEN_1046 : shotInteract_3; // @[Conditional.scala 39:67]
  wire  _GEN_1504 = _T_887 ? _GEN_1045 : shotPop_3; // @[Conditional.scala 39:67]
  wire  _GEN_1506 = _T_887 ? _GEN_1049 : spriteVisibleReg_6; // @[Conditional.scala 39:67]
  wire  _GEN_1507 = _T_887 ? _GEN_1052 : shotInteract_4; // @[Conditional.scala 39:67]
  wire  _GEN_1508 = _T_887 ? _GEN_1051 : shotPop_4; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_1517 = _T_887 ? _GEN_1059 : 2'h2; // @[Conditional.scala 39:67]
  wire  _GEN_1572 = _T_887 ? show : _GEN_1352; // @[Conditional.scala 39:67]
  wire  _GEN_1583 = _T_887 ? shipInteract : _GEN_1363; // @[Conditional.scala 39:67]
  wire  _GEN_1647 = _T_887 ? spriteVisibleReg_26 : _GEN_1427; // @[Conditional.scala 39:67]
  wire  _GEN_1650 = _T_887 ? spriteVisibleReg_30 : _GEN_1430; // @[Conditional.scala 39:67]
  wire  _GEN_1653 = _T_887 ? spriteVisibleReg_27 : _GEN_1433; // @[Conditional.scala 39:67]
  wire  _GEN_1656 = _T_887 ? spriteVisibleReg_31 : _GEN_1436; // @[Conditional.scala 39:67]
  wire  _GEN_1659 = _T_887 ? spriteVisibleReg_28 : _GEN_1439; // @[Conditional.scala 39:67]
  wire  _GEN_1662 = _T_887 ? spriteVisibleReg_32 : _GEN_1442; // @[Conditional.scala 39:67]
  wire  _GEN_1665 = _T_887 ? spriteVisibleReg_29 : _GEN_1445; // @[Conditional.scala 39:67]
  wire  _GEN_1668 = _T_887 ? spriteVisibleReg_33 : _GEN_1448; // @[Conditional.scala 39:67]
  wire  _GEN_1671 = _T_887 ? spriteVisibleReg_72 : _GEN_1451; // @[Conditional.scala 39:67]
  wire  _GEN_1672 = _T_887 ? spriteVisibleReg_66 : _GEN_1452; // @[Conditional.scala 39:67]
  wire  _GEN_1673 = _T_887 ? spriteVisibleReg_57 : _GEN_1453; // @[Conditional.scala 39:67]
  wire  _GEN_1674 = _T_887 ? spriteVisibleReg_61 : _GEN_1454; // @[Conditional.scala 39:67]
  wire  _GEN_1675 = _T_887 ? spriteVisibleReg_71 : _GEN_1455; // @[Conditional.scala 39:67]
  wire  _GEN_1676 = _T_887 ? spriteVisibleReg_65 : _GEN_1456; // @[Conditional.scala 39:67]
  wire  _GEN_1677 = _T_887 ? spriteVisibleReg_56 : _GEN_1457; // @[Conditional.scala 39:67]
  wire  _GEN_1678 = _T_887 ? spriteVisibleReg_62 : _GEN_1458; // @[Conditional.scala 39:67]
  wire  _GEN_1679 = _T_887 ? spriteVisibleReg_70 : _GEN_1459; // @[Conditional.scala 39:67]
  wire  _GEN_1680 = _T_887 ? spriteVisibleReg_64 : _GEN_1460; // @[Conditional.scala 39:67]
  wire  _GEN_1681 = _T_887 ? spriteVisibleReg_55 : _GEN_1461; // @[Conditional.scala 39:67]
  wire  _GEN_1682 = _T_887 ? spriteVisibleReg_63 : _GEN_1462; // @[Conditional.scala 39:67]
  wire  _GEN_1683 = _T_887 ? spriteVisibleReg_44 : _GEN_1463; // @[Conditional.scala 39:67]
  wire  _GEN_1686 = _T_887 ? spriteVisibleReg_45 : _GEN_1466; // @[Conditional.scala 39:67]
  wire  _GEN_1689 = _T_887 ? spriteVisibleReg_46 : _GEN_1469; // @[Conditional.scala 39:67]
  wire  _GEN_1692 = _T_887 ? spriteVisibleReg_47 : _GEN_1472; // @[Conditional.scala 39:67]
  wire  _GEN_1695 = _T_887 ? spriteVisibleReg_48 : _GEN_1475; // @[Conditional.scala 39:67]
  wire  _GEN_1698 = _T_887 ? spriteVisibleReg_49 : _GEN_1478; // @[Conditional.scala 39:67]
  wire  _GEN_1701 = _T_887 ? spriteVisibleReg_50 : _GEN_1481; // @[Conditional.scala 39:67]
  wire  _GEN_1704 = _T_887 ? spriteVisibleReg_51 : _GEN_1484; // @[Conditional.scala 39:67]
  wire  _GEN_1707 = _T_887 ? 1'h0 : _GEN_1488; // @[Conditional.scala 39:67]
  wire  _GEN_1712 = _T_863 ? spriteVisibleReg_2 : _GEN_1490; // @[Conditional.scala 39:67]
  wire  _GEN_1713 = _T_863 ? shotInteract_0 : _GEN_1491; // @[Conditional.scala 39:67]
  wire  _GEN_1714 = _T_863 ? shotPop_0 : _GEN_1492; // @[Conditional.scala 39:67]
  wire  _GEN_1716 = _T_863 ? spriteVisibleReg_3 : _GEN_1494; // @[Conditional.scala 39:67]
  wire  _GEN_1717 = _T_863 ? shotInteract_1 : _GEN_1495; // @[Conditional.scala 39:67]
  wire  _GEN_1718 = _T_863 ? shotPop_1 : _GEN_1496; // @[Conditional.scala 39:67]
  wire  _GEN_1720 = _T_863 ? spriteVisibleReg_4 : _GEN_1498; // @[Conditional.scala 39:67]
  wire  _GEN_1721 = _T_863 ? shotInteract_2 : _GEN_1499; // @[Conditional.scala 39:67]
  wire  _GEN_1722 = _T_863 ? shotPop_2 : _GEN_1500; // @[Conditional.scala 39:67]
  wire  _GEN_1724 = _T_863 ? spriteVisibleReg_5 : _GEN_1502; // @[Conditional.scala 39:67]
  wire  _GEN_1725 = _T_863 ? shotInteract_3 : _GEN_1503; // @[Conditional.scala 39:67]
  wire  _GEN_1726 = _T_863 ? shotPop_3 : _GEN_1504; // @[Conditional.scala 39:67]
  wire  _GEN_1728 = _T_863 ? spriteVisibleReg_6 : _GEN_1506; // @[Conditional.scala 39:67]
  wire  _GEN_1729 = _T_863 ? shotInteract_4 : _GEN_1507; // @[Conditional.scala 39:67]
  wire  _GEN_1730 = _T_863 ? shotPop_4 : _GEN_1508; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_1739 = _T_863 ? 2'h2 : _GEN_1517; // @[Conditional.scala 39:67]
  wire  _GEN_1793 = _T_863 ? show : _GEN_1572; // @[Conditional.scala 39:67]
  wire  _GEN_1802 = _T_863 ? shipInteract : _GEN_1583; // @[Conditional.scala 39:67]
  wire  _GEN_1866 = _T_863 ? spriteVisibleReg_26 : _GEN_1647; // @[Conditional.scala 39:67]
  wire  _GEN_1869 = _T_863 ? spriteVisibleReg_30 : _GEN_1650; // @[Conditional.scala 39:67]
  wire  _GEN_1872 = _T_863 ? spriteVisibleReg_27 : _GEN_1653; // @[Conditional.scala 39:67]
  wire  _GEN_1875 = _T_863 ? spriteVisibleReg_31 : _GEN_1656; // @[Conditional.scala 39:67]
  wire  _GEN_1878 = _T_863 ? spriteVisibleReg_28 : _GEN_1659; // @[Conditional.scala 39:67]
  wire  _GEN_1881 = _T_863 ? spriteVisibleReg_32 : _GEN_1662; // @[Conditional.scala 39:67]
  wire  _GEN_1884 = _T_863 ? spriteVisibleReg_29 : _GEN_1665; // @[Conditional.scala 39:67]
  wire  _GEN_1887 = _T_863 ? spriteVisibleReg_33 : _GEN_1668; // @[Conditional.scala 39:67]
  wire  _GEN_1890 = _T_863 ? spriteVisibleReg_72 : _GEN_1671; // @[Conditional.scala 39:67]
  wire  _GEN_1891 = _T_863 ? spriteVisibleReg_66 : _GEN_1672; // @[Conditional.scala 39:67]
  wire  _GEN_1892 = _T_863 ? spriteVisibleReg_57 : _GEN_1673; // @[Conditional.scala 39:67]
  wire  _GEN_1893 = _T_863 ? spriteVisibleReg_61 : _GEN_1674; // @[Conditional.scala 39:67]
  wire  _GEN_1894 = _T_863 ? spriteVisibleReg_71 : _GEN_1675; // @[Conditional.scala 39:67]
  wire  _GEN_1895 = _T_863 ? spriteVisibleReg_65 : _GEN_1676; // @[Conditional.scala 39:67]
  wire  _GEN_1896 = _T_863 ? spriteVisibleReg_56 : _GEN_1677; // @[Conditional.scala 39:67]
  wire  _GEN_1897 = _T_863 ? spriteVisibleReg_62 : _GEN_1678; // @[Conditional.scala 39:67]
  wire  _GEN_1898 = _T_863 ? spriteVisibleReg_70 : _GEN_1679; // @[Conditional.scala 39:67]
  wire  _GEN_1899 = _T_863 ? spriteVisibleReg_64 : _GEN_1680; // @[Conditional.scala 39:67]
  wire  _GEN_1900 = _T_863 ? spriteVisibleReg_55 : _GEN_1681; // @[Conditional.scala 39:67]
  wire  _GEN_1901 = _T_863 ? spriteVisibleReg_63 : _GEN_1682; // @[Conditional.scala 39:67]
  wire  _GEN_1902 = _T_863 ? spriteVisibleReg_44 : _GEN_1683; // @[Conditional.scala 39:67]
  wire  _GEN_1905 = _T_863 ? spriteVisibleReg_45 : _GEN_1686; // @[Conditional.scala 39:67]
  wire  _GEN_1908 = _T_863 ? spriteVisibleReg_46 : _GEN_1689; // @[Conditional.scala 39:67]
  wire  _GEN_1911 = _T_863 ? spriteVisibleReg_47 : _GEN_1692; // @[Conditional.scala 39:67]
  wire  _GEN_1914 = _T_863 ? spriteVisibleReg_48 : _GEN_1695; // @[Conditional.scala 39:67]
  wire  _GEN_1917 = _T_863 ? spriteVisibleReg_49 : _GEN_1698; // @[Conditional.scala 39:67]
  wire  _GEN_1920 = _T_863 ? spriteVisibleReg_50 : _GEN_1701; // @[Conditional.scala 39:67]
  wire  _GEN_1923 = _T_863 ? spriteVisibleReg_51 : _GEN_1704; // @[Conditional.scala 39:67]
  wire  _GEN_1926 = _T_863 ? 1'h0 : _GEN_1707; // @[Conditional.scala 39:67]
  wire  _GEN_1931 = _T_706 ? _GEN_836 : _GEN_1713; // @[Conditional.scala 39:67]
  wire  _GEN_1932 = _T_706 ? _GEN_837 : _GEN_1714; // @[Conditional.scala 39:67]
  wire  _GEN_1933 = _T_706 ? _GEN_838 : _GEN_1712; // @[Conditional.scala 39:67]
  wire  _GEN_1934 = _T_706 ? _GEN_841 : _GEN_1717; // @[Conditional.scala 39:67]
  wire  _GEN_1935 = _T_706 ? _GEN_842 : _GEN_1718; // @[Conditional.scala 39:67]
  wire  _GEN_1936 = _T_706 ? _GEN_843 : _GEN_1716; // @[Conditional.scala 39:67]
  wire  _GEN_1937 = _T_706 ? _GEN_846 : _GEN_1721; // @[Conditional.scala 39:67]
  wire  _GEN_1938 = _T_706 ? _GEN_847 : _GEN_1722; // @[Conditional.scala 39:67]
  wire  _GEN_1939 = _T_706 ? _GEN_848 : _GEN_1720; // @[Conditional.scala 39:67]
  wire  _GEN_1940 = _T_706 ? _GEN_851 : _GEN_1725; // @[Conditional.scala 39:67]
  wire  _GEN_1941 = _T_706 ? _GEN_852 : _GEN_1726; // @[Conditional.scala 39:67]
  wire  _GEN_1942 = _T_706 ? _GEN_853 : _GEN_1724; // @[Conditional.scala 39:67]
  wire  _GEN_1943 = _T_706 ? _GEN_856 : _GEN_1729; // @[Conditional.scala 39:67]
  wire  _GEN_1944 = _T_706 ? _GEN_857 : _GEN_1730; // @[Conditional.scala 39:67]
  wire  _GEN_1945 = _T_706 ? _GEN_858 : _GEN_1728; // @[Conditional.scala 39:67]
  wire  _GEN_1966 = _T_706 ? _GEN_825 : planetUp; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_1990 = _T_706 ? 2'h2 : _GEN_1739; // @[Conditional.scala 39:67]
  wire  _GEN_2030 = _T_706 ? show : _GEN_1793; // @[Conditional.scala 39:67]
  wire  _GEN_2039 = _T_706 ? shipInteract : _GEN_1802; // @[Conditional.scala 39:67]
  wire  _GEN_2102 = _T_706 ? spriteVisibleReg_26 : _GEN_1866; // @[Conditional.scala 39:67]
  wire  _GEN_2105 = _T_706 ? spriteVisibleReg_30 : _GEN_1869; // @[Conditional.scala 39:67]
  wire  _GEN_2108 = _T_706 ? spriteVisibleReg_27 : _GEN_1872; // @[Conditional.scala 39:67]
  wire  _GEN_2111 = _T_706 ? spriteVisibleReg_31 : _GEN_1875; // @[Conditional.scala 39:67]
  wire  _GEN_2114 = _T_706 ? spriteVisibleReg_28 : _GEN_1878; // @[Conditional.scala 39:67]
  wire  _GEN_2117 = _T_706 ? spriteVisibleReg_32 : _GEN_1881; // @[Conditional.scala 39:67]
  wire  _GEN_2120 = _T_706 ? spriteVisibleReg_29 : _GEN_1884; // @[Conditional.scala 39:67]
  wire  _GEN_2123 = _T_706 ? spriteVisibleReg_33 : _GEN_1887; // @[Conditional.scala 39:67]
  wire  _GEN_2126 = _T_706 ? spriteVisibleReg_72 : _GEN_1890; // @[Conditional.scala 39:67]
  wire  _GEN_2127 = _T_706 ? spriteVisibleReg_66 : _GEN_1891; // @[Conditional.scala 39:67]
  wire  _GEN_2128 = _T_706 ? spriteVisibleReg_57 : _GEN_1892; // @[Conditional.scala 39:67]
  wire  _GEN_2129 = _T_706 ? spriteVisibleReg_61 : _GEN_1893; // @[Conditional.scala 39:67]
  wire  _GEN_2130 = _T_706 ? spriteVisibleReg_71 : _GEN_1894; // @[Conditional.scala 39:67]
  wire  _GEN_2131 = _T_706 ? spriteVisibleReg_65 : _GEN_1895; // @[Conditional.scala 39:67]
  wire  _GEN_2132 = _T_706 ? spriteVisibleReg_56 : _GEN_1896; // @[Conditional.scala 39:67]
  wire  _GEN_2133 = _T_706 ? spriteVisibleReg_62 : _GEN_1897; // @[Conditional.scala 39:67]
  wire  _GEN_2134 = _T_706 ? spriteVisibleReg_70 : _GEN_1898; // @[Conditional.scala 39:67]
  wire  _GEN_2135 = _T_706 ? spriteVisibleReg_64 : _GEN_1899; // @[Conditional.scala 39:67]
  wire  _GEN_2136 = _T_706 ? spriteVisibleReg_55 : _GEN_1900; // @[Conditional.scala 39:67]
  wire  _GEN_2137 = _T_706 ? spriteVisibleReg_63 : _GEN_1901; // @[Conditional.scala 39:67]
  wire  _GEN_2138 = _T_706 ? spriteVisibleReg_44 : _GEN_1902; // @[Conditional.scala 39:67]
  wire  _GEN_2141 = _T_706 ? spriteVisibleReg_45 : _GEN_1905; // @[Conditional.scala 39:67]
  wire  _GEN_2144 = _T_706 ? spriteVisibleReg_46 : _GEN_1908; // @[Conditional.scala 39:67]
  wire  _GEN_2147 = _T_706 ? spriteVisibleReg_47 : _GEN_1911; // @[Conditional.scala 39:67]
  wire  _GEN_2150 = _T_706 ? spriteVisibleReg_48 : _GEN_1914; // @[Conditional.scala 39:67]
  wire  _GEN_2153 = _T_706 ? spriteVisibleReg_49 : _GEN_1917; // @[Conditional.scala 39:67]
  wire  _GEN_2156 = _T_706 ? spriteVisibleReg_50 : _GEN_1920; // @[Conditional.scala 39:67]
  wire  _GEN_2159 = _T_706 ? spriteVisibleReg_51 : _GEN_1923; // @[Conditional.scala 39:67]
  wire  _GEN_2162 = _T_706 ? 1'h0 : _GEN_1926; // @[Conditional.scala 39:67]
  wire  _GEN_2167 = _T_685 ? _GEN_593 : _GEN_1931; // @[Conditional.scala 39:67]
  wire  _GEN_2168 = _T_685 ? _GEN_594 : _GEN_1932; // @[Conditional.scala 39:67]
  wire  _GEN_2169 = _T_685 ? _GEN_595 : _GEN_1933; // @[Conditional.scala 39:67]
  wire  _GEN_2170 = _T_685 ? _GEN_596 : _GEN_1934; // @[Conditional.scala 39:67]
  wire  _GEN_2171 = _T_685 ? _GEN_597 : _GEN_1935; // @[Conditional.scala 39:67]
  wire  _GEN_2172 = _T_685 ? _GEN_598 : _GEN_1936; // @[Conditional.scala 39:67]
  wire  _GEN_2173 = _T_685 ? _GEN_599 : _GEN_1937; // @[Conditional.scala 39:67]
  wire  _GEN_2174 = _T_685 ? _GEN_600 : _GEN_1938; // @[Conditional.scala 39:67]
  wire  _GEN_2175 = _T_685 ? _GEN_601 : _GEN_1939; // @[Conditional.scala 39:67]
  wire  _GEN_2181 = _T_685 ? shotInteract_3 : _GEN_1940; // @[Conditional.scala 39:67]
  wire  _GEN_2182 = _T_685 ? shotPop_3 : _GEN_1941; // @[Conditional.scala 39:67]
  wire  _GEN_2183 = _T_685 ? spriteVisibleReg_5 : _GEN_1942; // @[Conditional.scala 39:67]
  wire  _GEN_2184 = _T_685 ? shotInteract_4 : _GEN_1943; // @[Conditional.scala 39:67]
  wire  _GEN_2185 = _T_685 ? shotPop_4 : _GEN_1944; // @[Conditional.scala 39:67]
  wire  _GEN_2186 = _T_685 ? spriteVisibleReg_6 : _GEN_1945; // @[Conditional.scala 39:67]
  wire  _GEN_2203 = _T_685 ? planetUp : _GEN_1966; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2226 = _T_685 ? 2'h2 : _GEN_1990; // @[Conditional.scala 39:67]
  wire  _GEN_2266 = _T_685 ? show : _GEN_2030; // @[Conditional.scala 39:67]
  wire  _GEN_2275 = _T_685 ? shipInteract : _GEN_2039; // @[Conditional.scala 39:67]
  wire  _GEN_2338 = _T_685 ? spriteVisibleReg_26 : _GEN_2102; // @[Conditional.scala 39:67]
  wire  _GEN_2341 = _T_685 ? spriteVisibleReg_30 : _GEN_2105; // @[Conditional.scala 39:67]
  wire  _GEN_2344 = _T_685 ? spriteVisibleReg_27 : _GEN_2108; // @[Conditional.scala 39:67]
  wire  _GEN_2347 = _T_685 ? spriteVisibleReg_31 : _GEN_2111; // @[Conditional.scala 39:67]
  wire  _GEN_2350 = _T_685 ? spriteVisibleReg_28 : _GEN_2114; // @[Conditional.scala 39:67]
  wire  _GEN_2353 = _T_685 ? spriteVisibleReg_32 : _GEN_2117; // @[Conditional.scala 39:67]
  wire  _GEN_2356 = _T_685 ? spriteVisibleReg_29 : _GEN_2120; // @[Conditional.scala 39:67]
  wire  _GEN_2359 = _T_685 ? spriteVisibleReg_33 : _GEN_2123; // @[Conditional.scala 39:67]
  wire  _GEN_2362 = _T_685 ? spriteVisibleReg_72 : _GEN_2126; // @[Conditional.scala 39:67]
  wire  _GEN_2363 = _T_685 ? spriteVisibleReg_66 : _GEN_2127; // @[Conditional.scala 39:67]
  wire  _GEN_2364 = _T_685 ? spriteVisibleReg_57 : _GEN_2128; // @[Conditional.scala 39:67]
  wire  _GEN_2365 = _T_685 ? spriteVisibleReg_61 : _GEN_2129; // @[Conditional.scala 39:67]
  wire  _GEN_2366 = _T_685 ? spriteVisibleReg_71 : _GEN_2130; // @[Conditional.scala 39:67]
  wire  _GEN_2367 = _T_685 ? spriteVisibleReg_65 : _GEN_2131; // @[Conditional.scala 39:67]
  wire  _GEN_2368 = _T_685 ? spriteVisibleReg_56 : _GEN_2132; // @[Conditional.scala 39:67]
  wire  _GEN_2369 = _T_685 ? spriteVisibleReg_62 : _GEN_2133; // @[Conditional.scala 39:67]
  wire  _GEN_2370 = _T_685 ? spriteVisibleReg_70 : _GEN_2134; // @[Conditional.scala 39:67]
  wire  _GEN_2371 = _T_685 ? spriteVisibleReg_64 : _GEN_2135; // @[Conditional.scala 39:67]
  wire  _GEN_2372 = _T_685 ? spriteVisibleReg_55 : _GEN_2136; // @[Conditional.scala 39:67]
  wire  _GEN_2373 = _T_685 ? spriteVisibleReg_63 : _GEN_2137; // @[Conditional.scala 39:67]
  wire  _GEN_2374 = _T_685 ? spriteVisibleReg_44 : _GEN_2138; // @[Conditional.scala 39:67]
  wire  _GEN_2377 = _T_685 ? spriteVisibleReg_45 : _GEN_2141; // @[Conditional.scala 39:67]
  wire  _GEN_2380 = _T_685 ? spriteVisibleReg_46 : _GEN_2144; // @[Conditional.scala 39:67]
  wire  _GEN_2383 = _T_685 ? spriteVisibleReg_47 : _GEN_2147; // @[Conditional.scala 39:67]
  wire  _GEN_2386 = _T_685 ? spriteVisibleReg_48 : _GEN_2150; // @[Conditional.scala 39:67]
  wire  _GEN_2389 = _T_685 ? spriteVisibleReg_49 : _GEN_2153; // @[Conditional.scala 39:67]
  wire  _GEN_2392 = _T_685 ? spriteVisibleReg_50 : _GEN_2156; // @[Conditional.scala 39:67]
  wire  _GEN_2395 = _T_685 ? spriteVisibleReg_51 : _GEN_2159; // @[Conditional.scala 39:67]
  wire  _GEN_2398 = _T_685 ? 1'h0 : _GEN_2162; // @[Conditional.scala 39:67]
  wire  _GEN_2403 = _T_628 ? _GEN_547 : _GEN_2167; // @[Conditional.scala 39:67]
  wire  _GEN_2404 = _T_628 ? _GEN_548 : _GEN_2168; // @[Conditional.scala 39:67]
  wire  _GEN_2405 = _T_628 ? _GEN_549 : _GEN_2169; // @[Conditional.scala 39:67]
  wire  _GEN_2406 = _T_628 ? _GEN_555 : _GEN_2170; // @[Conditional.scala 39:67]
  wire  _GEN_2407 = _T_628 ? _GEN_556 : _GEN_2171; // @[Conditional.scala 39:67]
  wire  _GEN_2408 = _T_628 ? _GEN_557 : _GEN_2172; // @[Conditional.scala 39:67]
  wire  _GEN_2409 = _T_628 ? _GEN_563 : _GEN_2173; // @[Conditional.scala 39:67]
  wire  _GEN_2410 = _T_628 ? _GEN_564 : _GEN_2174; // @[Conditional.scala 39:67]
  wire  _GEN_2411 = _T_628 ? _GEN_565 : _GEN_2175; // @[Conditional.scala 39:67]
  wire  _GEN_2412 = _T_628 ? _GEN_571 : _GEN_2181; // @[Conditional.scala 39:67]
  wire  _GEN_2413 = _T_628 ? _GEN_572 : _GEN_2182; // @[Conditional.scala 39:67]
  wire  _GEN_2414 = _T_628 ? _GEN_573 : _GEN_2183; // @[Conditional.scala 39:67]
  wire  _GEN_2415 = _T_628 ? _GEN_579 : _GEN_2184; // @[Conditional.scala 39:67]
  wire  _GEN_2416 = _T_628 ? _GEN_580 : _GEN_2185; // @[Conditional.scala 39:67]
  wire  _GEN_2417 = _T_628 ? _GEN_581 : _GEN_2186; // @[Conditional.scala 39:67]
  wire  _GEN_2451 = _T_628 ? planetUp : _GEN_2203; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2472 = _T_628 ? 2'h2 : _GEN_2226; // @[Conditional.scala 39:67]
  wire  _GEN_2508 = _T_628 ? show : _GEN_2266; // @[Conditional.scala 39:67]
  wire  _GEN_2517 = _T_628 ? shipInteract : _GEN_2275; // @[Conditional.scala 39:67]
  wire  _GEN_2580 = _T_628 ? spriteVisibleReg_26 : _GEN_2338; // @[Conditional.scala 39:67]
  wire  _GEN_2583 = _T_628 ? spriteVisibleReg_30 : _GEN_2341; // @[Conditional.scala 39:67]
  wire  _GEN_2586 = _T_628 ? spriteVisibleReg_27 : _GEN_2344; // @[Conditional.scala 39:67]
  wire  _GEN_2589 = _T_628 ? spriteVisibleReg_31 : _GEN_2347; // @[Conditional.scala 39:67]
  wire  _GEN_2592 = _T_628 ? spriteVisibleReg_28 : _GEN_2350; // @[Conditional.scala 39:67]
  wire  _GEN_2595 = _T_628 ? spriteVisibleReg_32 : _GEN_2353; // @[Conditional.scala 39:67]
  wire  _GEN_2598 = _T_628 ? spriteVisibleReg_29 : _GEN_2356; // @[Conditional.scala 39:67]
  wire  _GEN_2601 = _T_628 ? spriteVisibleReg_33 : _GEN_2359; // @[Conditional.scala 39:67]
  wire  _GEN_2604 = _T_628 ? spriteVisibleReg_72 : _GEN_2362; // @[Conditional.scala 39:67]
  wire  _GEN_2605 = _T_628 ? spriteVisibleReg_66 : _GEN_2363; // @[Conditional.scala 39:67]
  wire  _GEN_2606 = _T_628 ? spriteVisibleReg_57 : _GEN_2364; // @[Conditional.scala 39:67]
  wire  _GEN_2607 = _T_628 ? spriteVisibleReg_61 : _GEN_2365; // @[Conditional.scala 39:67]
  wire  _GEN_2608 = _T_628 ? spriteVisibleReg_71 : _GEN_2366; // @[Conditional.scala 39:67]
  wire  _GEN_2609 = _T_628 ? spriteVisibleReg_65 : _GEN_2367; // @[Conditional.scala 39:67]
  wire  _GEN_2610 = _T_628 ? spriteVisibleReg_56 : _GEN_2368; // @[Conditional.scala 39:67]
  wire  _GEN_2611 = _T_628 ? spriteVisibleReg_62 : _GEN_2369; // @[Conditional.scala 39:67]
  wire  _GEN_2612 = _T_628 ? spriteVisibleReg_70 : _GEN_2370; // @[Conditional.scala 39:67]
  wire  _GEN_2613 = _T_628 ? spriteVisibleReg_64 : _GEN_2371; // @[Conditional.scala 39:67]
  wire  _GEN_2614 = _T_628 ? spriteVisibleReg_55 : _GEN_2372; // @[Conditional.scala 39:67]
  wire  _GEN_2615 = _T_628 ? spriteVisibleReg_63 : _GEN_2373; // @[Conditional.scala 39:67]
  wire  _GEN_2616 = _T_628 ? spriteVisibleReg_44 : _GEN_2374; // @[Conditional.scala 39:67]
  wire  _GEN_2619 = _T_628 ? spriteVisibleReg_45 : _GEN_2377; // @[Conditional.scala 39:67]
  wire  _GEN_2622 = _T_628 ? spriteVisibleReg_46 : _GEN_2380; // @[Conditional.scala 39:67]
  wire  _GEN_2625 = _T_628 ? spriteVisibleReg_47 : _GEN_2383; // @[Conditional.scala 39:67]
  wire  _GEN_2628 = _T_628 ? spriteVisibleReg_48 : _GEN_2386; // @[Conditional.scala 39:67]
  wire  _GEN_2631 = _T_628 ? spriteVisibleReg_49 : _GEN_2389; // @[Conditional.scala 39:67]
  wire  _GEN_2634 = _T_628 ? spriteVisibleReg_50 : _GEN_2392; // @[Conditional.scala 39:67]
  wire  _GEN_2637 = _T_628 ? spriteVisibleReg_51 : _GEN_2395; // @[Conditional.scala 39:67]
  wire  _GEN_2640 = _T_628 ? 1'h0 : _GEN_2398; // @[Conditional.scala 39:67]
  wire  _GEN_2645 = _T_571 ? _GEN_397 : _GEN_2403; // @[Conditional.scala 39:67]
  wire  _GEN_2646 = _T_571 ? _GEN_398 : _GEN_2404; // @[Conditional.scala 39:67]
  wire  _GEN_2647 = _T_571 ? _GEN_399 : _GEN_2405; // @[Conditional.scala 39:67]
  wire  _GEN_2648 = _T_571 ? _GEN_405 : _GEN_2406; // @[Conditional.scala 39:67]
  wire  _GEN_2649 = _T_571 ? _GEN_406 : _GEN_2407; // @[Conditional.scala 39:67]
  wire  _GEN_2650 = _T_571 ? _GEN_407 : _GEN_2408; // @[Conditional.scala 39:67]
  wire  _GEN_2651 = _T_571 ? _GEN_413 : _GEN_2409; // @[Conditional.scala 39:67]
  wire  _GEN_2652 = _T_571 ? _GEN_414 : _GEN_2410; // @[Conditional.scala 39:67]
  wire  _GEN_2653 = _T_571 ? _GEN_415 : _GEN_2411; // @[Conditional.scala 39:67]
  wire  _GEN_2654 = _T_571 ? _GEN_421 : _GEN_2412; // @[Conditional.scala 39:67]
  wire  _GEN_2655 = _T_571 ? _GEN_422 : _GEN_2413; // @[Conditional.scala 39:67]
  wire  _GEN_2656 = _T_571 ? _GEN_423 : _GEN_2414; // @[Conditional.scala 39:67]
  wire  _GEN_2657 = _T_571 ? _GEN_429 : _GEN_2415; // @[Conditional.scala 39:67]
  wire  _GEN_2658 = _T_571 ? _GEN_430 : _GEN_2416; // @[Conditional.scala 39:67]
  wire  _GEN_2659 = _T_571 ? _GEN_431 : _GEN_2417; // @[Conditional.scala 39:67]
  wire  _GEN_2697 = _T_571 ? planetUp : _GEN_2451; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2718 = _T_571 ? 2'h2 : _GEN_2472; // @[Conditional.scala 39:67]
  wire  _GEN_2752 = _T_571 ? show : _GEN_2508; // @[Conditional.scala 39:67]
  wire  _GEN_2761 = _T_571 ? shipInteract : _GEN_2517; // @[Conditional.scala 39:67]
  wire  _GEN_2824 = _T_571 ? spriteVisibleReg_26 : _GEN_2580; // @[Conditional.scala 39:67]
  wire  _GEN_2827 = _T_571 ? spriteVisibleReg_30 : _GEN_2583; // @[Conditional.scala 39:67]
  wire  _GEN_2830 = _T_571 ? spriteVisibleReg_27 : _GEN_2586; // @[Conditional.scala 39:67]
  wire  _GEN_2833 = _T_571 ? spriteVisibleReg_31 : _GEN_2589; // @[Conditional.scala 39:67]
  wire  _GEN_2836 = _T_571 ? spriteVisibleReg_28 : _GEN_2592; // @[Conditional.scala 39:67]
  wire  _GEN_2839 = _T_571 ? spriteVisibleReg_32 : _GEN_2595; // @[Conditional.scala 39:67]
  wire  _GEN_2842 = _T_571 ? spriteVisibleReg_29 : _GEN_2598; // @[Conditional.scala 39:67]
  wire  _GEN_2845 = _T_571 ? spriteVisibleReg_33 : _GEN_2601; // @[Conditional.scala 39:67]
  wire  _GEN_2848 = _T_571 ? spriteVisibleReg_72 : _GEN_2604; // @[Conditional.scala 39:67]
  wire  _GEN_2849 = _T_571 ? spriteVisibleReg_66 : _GEN_2605; // @[Conditional.scala 39:67]
  wire  _GEN_2850 = _T_571 ? spriteVisibleReg_57 : _GEN_2606; // @[Conditional.scala 39:67]
  wire  _GEN_2851 = _T_571 ? spriteVisibleReg_61 : _GEN_2607; // @[Conditional.scala 39:67]
  wire  _GEN_2852 = _T_571 ? spriteVisibleReg_71 : _GEN_2608; // @[Conditional.scala 39:67]
  wire  _GEN_2853 = _T_571 ? spriteVisibleReg_65 : _GEN_2609; // @[Conditional.scala 39:67]
  wire  _GEN_2854 = _T_571 ? spriteVisibleReg_56 : _GEN_2610; // @[Conditional.scala 39:67]
  wire  _GEN_2855 = _T_571 ? spriteVisibleReg_62 : _GEN_2611; // @[Conditional.scala 39:67]
  wire  _GEN_2856 = _T_571 ? spriteVisibleReg_70 : _GEN_2612; // @[Conditional.scala 39:67]
  wire  _GEN_2857 = _T_571 ? spriteVisibleReg_64 : _GEN_2613; // @[Conditional.scala 39:67]
  wire  _GEN_2858 = _T_571 ? spriteVisibleReg_55 : _GEN_2614; // @[Conditional.scala 39:67]
  wire  _GEN_2859 = _T_571 ? spriteVisibleReg_63 : _GEN_2615; // @[Conditional.scala 39:67]
  wire  _GEN_2860 = _T_571 ? spriteVisibleReg_44 : _GEN_2616; // @[Conditional.scala 39:67]
  wire  _GEN_2863 = _T_571 ? spriteVisibleReg_45 : _GEN_2619; // @[Conditional.scala 39:67]
  wire  _GEN_2866 = _T_571 ? spriteVisibleReg_46 : _GEN_2622; // @[Conditional.scala 39:67]
  wire  _GEN_2869 = _T_571 ? spriteVisibleReg_47 : _GEN_2625; // @[Conditional.scala 39:67]
  wire  _GEN_2872 = _T_571 ? spriteVisibleReg_48 : _GEN_2628; // @[Conditional.scala 39:67]
  wire  _GEN_2875 = _T_571 ? spriteVisibleReg_49 : _GEN_2631; // @[Conditional.scala 39:67]
  wire  _GEN_2878 = _T_571 ? spriteVisibleReg_50 : _GEN_2634; // @[Conditional.scala 39:67]
  wire  _GEN_2881 = _T_571 ? spriteVisibleReg_51 : _GEN_2637; // @[Conditional.scala 39:67]
  wire  _GEN_2884 = _T_571 ? 1'h0 : _GEN_2640; // @[Conditional.scala 39:67]
  wire  _GEN_2889 = _T_506 ? _GEN_259 : _GEN_2645; // @[Conditional.scala 39:67]
  wire  _GEN_2890 = _T_506 ? _GEN_260 : _GEN_2646; // @[Conditional.scala 39:67]
  wire  _GEN_2891 = _T_506 ? _GEN_261 : _GEN_2647; // @[Conditional.scala 39:67]
  wire  _GEN_2892 = _T_506 ? _GEN_262 : _GEN_2648; // @[Conditional.scala 39:67]
  wire  _GEN_2893 = _T_506 ? _GEN_263 : _GEN_2649; // @[Conditional.scala 39:67]
  wire  _GEN_2894 = _T_506 ? _GEN_264 : _GEN_2650; // @[Conditional.scala 39:67]
  wire  _GEN_2895 = _T_506 ? _GEN_265 : _GEN_2651; // @[Conditional.scala 39:67]
  wire  _GEN_2896 = _T_506 ? _GEN_266 : _GEN_2652; // @[Conditional.scala 39:67]
  wire  _GEN_2897 = _T_506 ? _GEN_267 : _GEN_2653; // @[Conditional.scala 39:67]
  wire  _GEN_2898 = _T_506 ? _GEN_268 : _GEN_2654; // @[Conditional.scala 39:67]
  wire  _GEN_2899 = _T_506 ? _GEN_269 : _GEN_2655; // @[Conditional.scala 39:67]
  wire  _GEN_2900 = _T_506 ? _GEN_270 : _GEN_2656; // @[Conditional.scala 39:67]
  wire  _GEN_2901 = _T_506 ? _GEN_271 : _GEN_2657; // @[Conditional.scala 39:67]
  wire  _GEN_2902 = _T_506 ? _GEN_272 : _GEN_2658; // @[Conditional.scala 39:67]
  wire  _GEN_2903 = _T_506 ? _GEN_273 : _GEN_2659; // @[Conditional.scala 39:67]
  wire  _GEN_2941 = _T_506 ? planetUp : _GEN_2697; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2962 = _T_506 ? 2'h2 : _GEN_2718; // @[Conditional.scala 39:67]
  wire  _GEN_2996 = _T_506 ? show : _GEN_2752; // @[Conditional.scala 39:67]
  wire  _GEN_3005 = _T_506 ? shipInteract : _GEN_2761; // @[Conditional.scala 39:67]
  wire  _GEN_3068 = _T_506 ? spriteVisibleReg_26 : _GEN_2824; // @[Conditional.scala 39:67]
  wire  _GEN_3071 = _T_506 ? spriteVisibleReg_30 : _GEN_2827; // @[Conditional.scala 39:67]
  wire  _GEN_3074 = _T_506 ? spriteVisibleReg_27 : _GEN_2830; // @[Conditional.scala 39:67]
  wire  _GEN_3077 = _T_506 ? spriteVisibleReg_31 : _GEN_2833; // @[Conditional.scala 39:67]
  wire  _GEN_3080 = _T_506 ? spriteVisibleReg_28 : _GEN_2836; // @[Conditional.scala 39:67]
  wire  _GEN_3083 = _T_506 ? spriteVisibleReg_32 : _GEN_2839; // @[Conditional.scala 39:67]
  wire  _GEN_3086 = _T_506 ? spriteVisibleReg_29 : _GEN_2842; // @[Conditional.scala 39:67]
  wire  _GEN_3089 = _T_506 ? spriteVisibleReg_33 : _GEN_2845; // @[Conditional.scala 39:67]
  wire  _GEN_3092 = _T_506 ? spriteVisibleReg_72 : _GEN_2848; // @[Conditional.scala 39:67]
  wire  _GEN_3093 = _T_506 ? spriteVisibleReg_66 : _GEN_2849; // @[Conditional.scala 39:67]
  wire  _GEN_3094 = _T_506 ? spriteVisibleReg_57 : _GEN_2850; // @[Conditional.scala 39:67]
  wire  _GEN_3095 = _T_506 ? spriteVisibleReg_61 : _GEN_2851; // @[Conditional.scala 39:67]
  wire  _GEN_3096 = _T_506 ? spriteVisibleReg_71 : _GEN_2852; // @[Conditional.scala 39:67]
  wire  _GEN_3097 = _T_506 ? spriteVisibleReg_65 : _GEN_2853; // @[Conditional.scala 39:67]
  wire  _GEN_3098 = _T_506 ? spriteVisibleReg_56 : _GEN_2854; // @[Conditional.scala 39:67]
  wire  _GEN_3099 = _T_506 ? spriteVisibleReg_62 : _GEN_2855; // @[Conditional.scala 39:67]
  wire  _GEN_3100 = _T_506 ? spriteVisibleReg_70 : _GEN_2856; // @[Conditional.scala 39:67]
  wire  _GEN_3101 = _T_506 ? spriteVisibleReg_64 : _GEN_2857; // @[Conditional.scala 39:67]
  wire  _GEN_3102 = _T_506 ? spriteVisibleReg_55 : _GEN_2858; // @[Conditional.scala 39:67]
  wire  _GEN_3103 = _T_506 ? spriteVisibleReg_63 : _GEN_2859; // @[Conditional.scala 39:67]
  wire  _GEN_3104 = _T_506 ? spriteVisibleReg_44 : _GEN_2860; // @[Conditional.scala 39:67]
  wire  _GEN_3107 = _T_506 ? spriteVisibleReg_45 : _GEN_2863; // @[Conditional.scala 39:67]
  wire  _GEN_3110 = _T_506 ? spriteVisibleReg_46 : _GEN_2866; // @[Conditional.scala 39:67]
  wire  _GEN_3113 = _T_506 ? spriteVisibleReg_47 : _GEN_2869; // @[Conditional.scala 39:67]
  wire  _GEN_3116 = _T_506 ? spriteVisibleReg_48 : _GEN_2872; // @[Conditional.scala 39:67]
  wire  _GEN_3119 = _T_506 ? spriteVisibleReg_49 : _GEN_2875; // @[Conditional.scala 39:67]
  wire  _GEN_3122 = _T_506 ? spriteVisibleReg_50 : _GEN_2878; // @[Conditional.scala 39:67]
  wire  _GEN_3125 = _T_506 ? spriteVisibleReg_51 : _GEN_2881; // @[Conditional.scala 39:67]
  wire  _GEN_3128 = _T_506 ? 1'h0 : _GEN_2884; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3129 = _T_487 ? _GEN_76 : 6'h0; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3130 = _T_487 ? _GEN_101 : 13'h0; // @[Conditional.scala 39:67]
  wire  _GEN_3131 = _T_487 & _T_409; // @[Conditional.scala 39:67]
  wire  _GEN_3138 = _T_487 ? shotInteract_0 : _GEN_2889; // @[Conditional.scala 39:67]
  wire  _GEN_3139 = _T_487 ? shotPop_0 : _GEN_2890; // @[Conditional.scala 39:67]
  wire  _GEN_3140 = _T_487 ? spriteVisibleReg_2 : _GEN_2891; // @[Conditional.scala 39:67]
  wire  _GEN_3141 = _T_487 ? shotInteract_1 : _GEN_2892; // @[Conditional.scala 39:67]
  wire  _GEN_3142 = _T_487 ? shotPop_1 : _GEN_2893; // @[Conditional.scala 39:67]
  wire  _GEN_3143 = _T_487 ? spriteVisibleReg_3 : _GEN_2894; // @[Conditional.scala 39:67]
  wire  _GEN_3144 = _T_487 ? shotInteract_2 : _GEN_2895; // @[Conditional.scala 39:67]
  wire  _GEN_3145 = _T_487 ? shotPop_2 : _GEN_2896; // @[Conditional.scala 39:67]
  wire  _GEN_3146 = _T_487 ? spriteVisibleReg_4 : _GEN_2897; // @[Conditional.scala 39:67]
  wire  _GEN_3147 = _T_487 ? shotInteract_3 : _GEN_2898; // @[Conditional.scala 39:67]
  wire  _GEN_3148 = _T_487 ? shotPop_3 : _GEN_2899; // @[Conditional.scala 39:67]
  wire  _GEN_3149 = _T_487 ? spriteVisibleReg_5 : _GEN_2900; // @[Conditional.scala 39:67]
  wire  _GEN_3150 = _T_487 ? shotInteract_4 : _GEN_2901; // @[Conditional.scala 39:67]
  wire  _GEN_3151 = _T_487 ? shotPop_4 : _GEN_2902; // @[Conditional.scala 39:67]
  wire  _GEN_3152 = _T_487 ? spriteVisibleReg_6 : _GEN_2903; // @[Conditional.scala 39:67]
  wire  _GEN_3189 = _T_487 ? planetUp : _GEN_2941; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3210 = _T_487 ? 2'h2 : _GEN_2962; // @[Conditional.scala 39:67]
  wire  _GEN_3244 = _T_487 ? show : _GEN_2996; // @[Conditional.scala 39:67]
  wire  _GEN_3253 = _T_487 ? shipInteract : _GEN_3005; // @[Conditional.scala 39:67]
  wire  _GEN_3316 = _T_487 ? spriteVisibleReg_26 : _GEN_3068; // @[Conditional.scala 39:67]
  wire  _GEN_3319 = _T_487 ? spriteVisibleReg_30 : _GEN_3071; // @[Conditional.scala 39:67]
  wire  _GEN_3322 = _T_487 ? spriteVisibleReg_27 : _GEN_3074; // @[Conditional.scala 39:67]
  wire  _GEN_3325 = _T_487 ? spriteVisibleReg_31 : _GEN_3077; // @[Conditional.scala 39:67]
  wire  _GEN_3328 = _T_487 ? spriteVisibleReg_28 : _GEN_3080; // @[Conditional.scala 39:67]
  wire  _GEN_3331 = _T_487 ? spriteVisibleReg_32 : _GEN_3083; // @[Conditional.scala 39:67]
  wire  _GEN_3334 = _T_487 ? spriteVisibleReg_29 : _GEN_3086; // @[Conditional.scala 39:67]
  wire  _GEN_3337 = _T_487 ? spriteVisibleReg_33 : _GEN_3089; // @[Conditional.scala 39:67]
  wire  _GEN_3340 = _T_487 ? spriteVisibleReg_72 : _GEN_3092; // @[Conditional.scala 39:67]
  wire  _GEN_3341 = _T_487 ? spriteVisibleReg_66 : _GEN_3093; // @[Conditional.scala 39:67]
  wire  _GEN_3342 = _T_487 ? spriteVisibleReg_57 : _GEN_3094; // @[Conditional.scala 39:67]
  wire  _GEN_3343 = _T_487 ? spriteVisibleReg_61 : _GEN_3095; // @[Conditional.scala 39:67]
  wire  _GEN_3344 = _T_487 ? spriteVisibleReg_71 : _GEN_3096; // @[Conditional.scala 39:67]
  wire  _GEN_3345 = _T_487 ? spriteVisibleReg_65 : _GEN_3097; // @[Conditional.scala 39:67]
  wire  _GEN_3346 = _T_487 ? spriteVisibleReg_56 : _GEN_3098; // @[Conditional.scala 39:67]
  wire  _GEN_3347 = _T_487 ? spriteVisibleReg_62 : _GEN_3099; // @[Conditional.scala 39:67]
  wire  _GEN_3348 = _T_487 ? spriteVisibleReg_70 : _GEN_3100; // @[Conditional.scala 39:67]
  wire  _GEN_3349 = _T_487 ? spriteVisibleReg_64 : _GEN_3101; // @[Conditional.scala 39:67]
  wire  _GEN_3350 = _T_487 ? spriteVisibleReg_55 : _GEN_3102; // @[Conditional.scala 39:67]
  wire  _GEN_3351 = _T_487 ? spriteVisibleReg_63 : _GEN_3103; // @[Conditional.scala 39:67]
  wire  _GEN_3352 = _T_487 ? spriteVisibleReg_44 : _GEN_3104; // @[Conditional.scala 39:67]
  wire  _GEN_3355 = _T_487 ? spriteVisibleReg_45 : _GEN_3107; // @[Conditional.scala 39:67]
  wire  _GEN_3358 = _T_487 ? spriteVisibleReg_46 : _GEN_3110; // @[Conditional.scala 39:67]
  wire  _GEN_3361 = _T_487 ? spriteVisibleReg_47 : _GEN_3113; // @[Conditional.scala 39:67]
  wire  _GEN_3364 = _T_487 ? spriteVisibleReg_48 : _GEN_3116; // @[Conditional.scala 39:67]
  wire  _GEN_3367 = _T_487 ? spriteVisibleReg_49 : _GEN_3119; // @[Conditional.scala 39:67]
  wire  _GEN_3370 = _T_487 ? spriteVisibleReg_50 : _GEN_3122; // @[Conditional.scala 39:67]
  wire  _GEN_3373 = _T_487 ? spriteVisibleReg_51 : _GEN_3125; // @[Conditional.scala 39:67]
  wire  _GEN_3376 = _T_487 ? 1'h0 : _GEN_3128; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3380 = _T_452 ? _GEN_93 : _GEN_3129; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3381 = _T_452 ? _GEN_94 : _GEN_3130; // @[Conditional.scala 39:67]
  wire  _GEN_3382 = _T_452 ? _GEN_95 : _GEN_3131; // @[Conditional.scala 39:67]
  wire  _GEN_3388 = _T_452 ? shotInteract_0 : _GEN_3138; // @[Conditional.scala 39:67]
  wire  _GEN_3389 = _T_452 ? shotPop_0 : _GEN_3139; // @[Conditional.scala 39:67]
  wire  _GEN_3390 = _T_452 ? spriteVisibleReg_2 : _GEN_3140; // @[Conditional.scala 39:67]
  wire  _GEN_3391 = _T_452 ? shotInteract_1 : _GEN_3141; // @[Conditional.scala 39:67]
  wire  _GEN_3392 = _T_452 ? shotPop_1 : _GEN_3142; // @[Conditional.scala 39:67]
  wire  _GEN_3393 = _T_452 ? spriteVisibleReg_3 : _GEN_3143; // @[Conditional.scala 39:67]
  wire  _GEN_3394 = _T_452 ? shotInteract_2 : _GEN_3144; // @[Conditional.scala 39:67]
  wire  _GEN_3395 = _T_452 ? shotPop_2 : _GEN_3145; // @[Conditional.scala 39:67]
  wire  _GEN_3396 = _T_452 ? spriteVisibleReg_4 : _GEN_3146; // @[Conditional.scala 39:67]
  wire  _GEN_3397 = _T_452 ? shotInteract_3 : _GEN_3147; // @[Conditional.scala 39:67]
  wire  _GEN_3398 = _T_452 ? shotPop_3 : _GEN_3148; // @[Conditional.scala 39:67]
  wire  _GEN_3399 = _T_452 ? spriteVisibleReg_5 : _GEN_3149; // @[Conditional.scala 39:67]
  wire  _GEN_3400 = _T_452 ? shotInteract_4 : _GEN_3150; // @[Conditional.scala 39:67]
  wire  _GEN_3401 = _T_452 ? shotPop_4 : _GEN_3151; // @[Conditional.scala 39:67]
  wire  _GEN_3402 = _T_452 ? spriteVisibleReg_6 : _GEN_3152; // @[Conditional.scala 39:67]
  wire  _GEN_3439 = _T_452 ? planetUp : _GEN_3189; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3460 = _T_452 ? 2'h2 : _GEN_3210; // @[Conditional.scala 39:67]
  wire  _GEN_3494 = _T_452 ? show : _GEN_3244; // @[Conditional.scala 39:67]
  wire  _GEN_3503 = _T_452 ? shipInteract : _GEN_3253; // @[Conditional.scala 39:67]
  wire  _GEN_3566 = _T_452 ? spriteVisibleReg_26 : _GEN_3316; // @[Conditional.scala 39:67]
  wire  _GEN_3569 = _T_452 ? spriteVisibleReg_30 : _GEN_3319; // @[Conditional.scala 39:67]
  wire  _GEN_3572 = _T_452 ? spriteVisibleReg_27 : _GEN_3322; // @[Conditional.scala 39:67]
  wire  _GEN_3575 = _T_452 ? spriteVisibleReg_31 : _GEN_3325; // @[Conditional.scala 39:67]
  wire  _GEN_3578 = _T_452 ? spriteVisibleReg_28 : _GEN_3328; // @[Conditional.scala 39:67]
  wire  _GEN_3581 = _T_452 ? spriteVisibleReg_32 : _GEN_3331; // @[Conditional.scala 39:67]
  wire  _GEN_3584 = _T_452 ? spriteVisibleReg_29 : _GEN_3334; // @[Conditional.scala 39:67]
  wire  _GEN_3587 = _T_452 ? spriteVisibleReg_33 : _GEN_3337; // @[Conditional.scala 39:67]
  wire  _GEN_3590 = _T_452 ? spriteVisibleReg_72 : _GEN_3340; // @[Conditional.scala 39:67]
  wire  _GEN_3591 = _T_452 ? spriteVisibleReg_66 : _GEN_3341; // @[Conditional.scala 39:67]
  wire  _GEN_3592 = _T_452 ? spriteVisibleReg_57 : _GEN_3342; // @[Conditional.scala 39:67]
  wire  _GEN_3593 = _T_452 ? spriteVisibleReg_61 : _GEN_3343; // @[Conditional.scala 39:67]
  wire  _GEN_3594 = _T_452 ? spriteVisibleReg_71 : _GEN_3344; // @[Conditional.scala 39:67]
  wire  _GEN_3595 = _T_452 ? spriteVisibleReg_65 : _GEN_3345; // @[Conditional.scala 39:67]
  wire  _GEN_3596 = _T_452 ? spriteVisibleReg_56 : _GEN_3346; // @[Conditional.scala 39:67]
  wire  _GEN_3597 = _T_452 ? spriteVisibleReg_62 : _GEN_3347; // @[Conditional.scala 39:67]
  wire  _GEN_3598 = _T_452 ? spriteVisibleReg_70 : _GEN_3348; // @[Conditional.scala 39:67]
  wire  _GEN_3599 = _T_452 ? spriteVisibleReg_64 : _GEN_3349; // @[Conditional.scala 39:67]
  wire  _GEN_3600 = _T_452 ? spriteVisibleReg_55 : _GEN_3350; // @[Conditional.scala 39:67]
  wire  _GEN_3601 = _T_452 ? spriteVisibleReg_63 : _GEN_3351; // @[Conditional.scala 39:67]
  wire  _GEN_3602 = _T_452 ? spriteVisibleReg_44 : _GEN_3352; // @[Conditional.scala 39:67]
  wire  _GEN_3605 = _T_452 ? spriteVisibleReg_45 : _GEN_3355; // @[Conditional.scala 39:67]
  wire  _GEN_3608 = _T_452 ? spriteVisibleReg_46 : _GEN_3358; // @[Conditional.scala 39:67]
  wire  _GEN_3611 = _T_452 ? spriteVisibleReg_47 : _GEN_3361; // @[Conditional.scala 39:67]
  wire  _GEN_3614 = _T_452 ? spriteVisibleReg_48 : _GEN_3364; // @[Conditional.scala 39:67]
  wire  _GEN_3617 = _T_452 ? spriteVisibleReg_49 : _GEN_3367; // @[Conditional.scala 39:67]
  wire  _GEN_3620 = _T_452 ? spriteVisibleReg_50 : _GEN_3370; // @[Conditional.scala 39:67]
  wire  _GEN_3623 = _T_452 ? spriteVisibleReg_51 : _GEN_3373; // @[Conditional.scala 39:67]
  wire  _GEN_3626 = _T_452 ? 1'h0 : _GEN_3376; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3630 = _T_405 ? _GEN_67 : _GEN_3380; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3631 = _T_405 ? _GEN_68 : _GEN_3381; // @[Conditional.scala 39:67]
  wire  _GEN_3632 = _T_405 ? _GEN_69 : _GEN_3382; // @[Conditional.scala 39:67]
  wire  _GEN_3639 = _T_405 ? shotInteract_0 : _GEN_3388; // @[Conditional.scala 39:67]
  wire  _GEN_3640 = _T_405 ? shotPop_0 : _GEN_3389; // @[Conditional.scala 39:67]
  wire  _GEN_3641 = _T_405 ? spriteVisibleReg_2 : _GEN_3390; // @[Conditional.scala 39:67]
  wire  _GEN_3642 = _T_405 ? shotInteract_1 : _GEN_3391; // @[Conditional.scala 39:67]
  wire  _GEN_3643 = _T_405 ? shotPop_1 : _GEN_3392; // @[Conditional.scala 39:67]
  wire  _GEN_3644 = _T_405 ? spriteVisibleReg_3 : _GEN_3393; // @[Conditional.scala 39:67]
  wire  _GEN_3645 = _T_405 ? shotInteract_2 : _GEN_3394; // @[Conditional.scala 39:67]
  wire  _GEN_3646 = _T_405 ? shotPop_2 : _GEN_3395; // @[Conditional.scala 39:67]
  wire  _GEN_3647 = _T_405 ? spriteVisibleReg_4 : _GEN_3396; // @[Conditional.scala 39:67]
  wire  _GEN_3648 = _T_405 ? shotInteract_3 : _GEN_3397; // @[Conditional.scala 39:67]
  wire  _GEN_3649 = _T_405 ? shotPop_3 : _GEN_3398; // @[Conditional.scala 39:67]
  wire  _GEN_3650 = _T_405 ? spriteVisibleReg_5 : _GEN_3399; // @[Conditional.scala 39:67]
  wire  _GEN_3651 = _T_405 ? shotInteract_4 : _GEN_3400; // @[Conditional.scala 39:67]
  wire  _GEN_3652 = _T_405 ? shotPop_4 : _GEN_3401; // @[Conditional.scala 39:67]
  wire  _GEN_3653 = _T_405 ? spriteVisibleReg_6 : _GEN_3402; // @[Conditional.scala 39:67]
  wire  _GEN_3690 = _T_405 ? planetUp : _GEN_3439; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3711 = _T_405 ? 2'h2 : _GEN_3460; // @[Conditional.scala 39:67]
  wire  _GEN_3744 = _T_405 ? show : _GEN_3494; // @[Conditional.scala 39:67]
  wire  _GEN_3753 = _T_405 ? shipInteract : _GEN_3503; // @[Conditional.scala 39:67]
  wire  _GEN_3816 = _T_405 ? spriteVisibleReg_26 : _GEN_3566; // @[Conditional.scala 39:67]
  wire  _GEN_3819 = _T_405 ? spriteVisibleReg_30 : _GEN_3569; // @[Conditional.scala 39:67]
  wire  _GEN_3822 = _T_405 ? spriteVisibleReg_27 : _GEN_3572; // @[Conditional.scala 39:67]
  wire  _GEN_3825 = _T_405 ? spriteVisibleReg_31 : _GEN_3575; // @[Conditional.scala 39:67]
  wire  _GEN_3828 = _T_405 ? spriteVisibleReg_28 : _GEN_3578; // @[Conditional.scala 39:67]
  wire  _GEN_3831 = _T_405 ? spriteVisibleReg_32 : _GEN_3581; // @[Conditional.scala 39:67]
  wire  _GEN_3834 = _T_405 ? spriteVisibleReg_29 : _GEN_3584; // @[Conditional.scala 39:67]
  wire  _GEN_3837 = _T_405 ? spriteVisibleReg_33 : _GEN_3587; // @[Conditional.scala 39:67]
  wire  _GEN_3840 = _T_405 ? spriteVisibleReg_72 : _GEN_3590; // @[Conditional.scala 39:67]
  wire  _GEN_3841 = _T_405 ? spriteVisibleReg_66 : _GEN_3591; // @[Conditional.scala 39:67]
  wire  _GEN_3842 = _T_405 ? spriteVisibleReg_57 : _GEN_3592; // @[Conditional.scala 39:67]
  wire  _GEN_3843 = _T_405 ? spriteVisibleReg_61 : _GEN_3593; // @[Conditional.scala 39:67]
  wire  _GEN_3844 = _T_405 ? spriteVisibleReg_71 : _GEN_3594; // @[Conditional.scala 39:67]
  wire  _GEN_3845 = _T_405 ? spriteVisibleReg_65 : _GEN_3595; // @[Conditional.scala 39:67]
  wire  _GEN_3846 = _T_405 ? spriteVisibleReg_56 : _GEN_3596; // @[Conditional.scala 39:67]
  wire  _GEN_3847 = _T_405 ? spriteVisibleReg_62 : _GEN_3597; // @[Conditional.scala 39:67]
  wire  _GEN_3848 = _T_405 ? spriteVisibleReg_70 : _GEN_3598; // @[Conditional.scala 39:67]
  wire  _GEN_3849 = _T_405 ? spriteVisibleReg_64 : _GEN_3599; // @[Conditional.scala 39:67]
  wire  _GEN_3850 = _T_405 ? spriteVisibleReg_55 : _GEN_3600; // @[Conditional.scala 39:67]
  wire  _GEN_3851 = _T_405 ? spriteVisibleReg_63 : _GEN_3601; // @[Conditional.scala 39:67]
  wire  _GEN_3852 = _T_405 ? spriteVisibleReg_44 : _GEN_3602; // @[Conditional.scala 39:67]
  wire  _GEN_3855 = _T_405 ? spriteVisibleReg_45 : _GEN_3605; // @[Conditional.scala 39:67]
  wire  _GEN_3858 = _T_405 ? spriteVisibleReg_46 : _GEN_3608; // @[Conditional.scala 39:67]
  wire  _GEN_3861 = _T_405 ? spriteVisibleReg_47 : _GEN_3611; // @[Conditional.scala 39:67]
  wire  _GEN_3864 = _T_405 ? spriteVisibleReg_48 : _GEN_3614; // @[Conditional.scala 39:67]
  wire  _GEN_3867 = _T_405 ? spriteVisibleReg_49 : _GEN_3617; // @[Conditional.scala 39:67]
  wire  _GEN_3870 = _T_405 ? spriteVisibleReg_50 : _GEN_3620; // @[Conditional.scala 39:67]
  wire  _GEN_3873 = _T_405 ? spriteVisibleReg_51 : _GEN_3623; // @[Conditional.scala 39:67]
  wire  _GEN_3876 = _T_405 ? 1'h0 : _GEN_3626; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3897 = _T_343 ? 6'h0 : _GEN_3630; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3898 = _T_343 ? 13'h0 : _GEN_3631; // @[Conditional.scala 39:67]
  wire  _GEN_3899 = _T_343 ? 1'h0 : _GEN_3632; // @[Conditional.scala 39:67]
  wire  _GEN_3905 = _T_343 ? shotInteract_0 : _GEN_3639; // @[Conditional.scala 39:67]
  wire  _GEN_3906 = _T_343 ? shotPop_0 : _GEN_3640; // @[Conditional.scala 39:67]
  wire  _GEN_3907 = _T_343 ? spriteVisibleReg_2 : _GEN_3641; // @[Conditional.scala 39:67]
  wire  _GEN_3908 = _T_343 ? shotInteract_1 : _GEN_3642; // @[Conditional.scala 39:67]
  wire  _GEN_3909 = _T_343 ? shotPop_1 : _GEN_3643; // @[Conditional.scala 39:67]
  wire  _GEN_3910 = _T_343 ? spriteVisibleReg_3 : _GEN_3644; // @[Conditional.scala 39:67]
  wire  _GEN_3911 = _T_343 ? shotInteract_2 : _GEN_3645; // @[Conditional.scala 39:67]
  wire  _GEN_3912 = _T_343 ? shotPop_2 : _GEN_3646; // @[Conditional.scala 39:67]
  wire  _GEN_3913 = _T_343 ? spriteVisibleReg_4 : _GEN_3647; // @[Conditional.scala 39:67]
  wire  _GEN_3914 = _T_343 ? shotInteract_3 : _GEN_3648; // @[Conditional.scala 39:67]
  wire  _GEN_3915 = _T_343 ? shotPop_3 : _GEN_3649; // @[Conditional.scala 39:67]
  wire  _GEN_3916 = _T_343 ? spriteVisibleReg_5 : _GEN_3650; // @[Conditional.scala 39:67]
  wire  _GEN_3917 = _T_343 ? shotInteract_4 : _GEN_3651; // @[Conditional.scala 39:67]
  wire  _GEN_3918 = _T_343 ? shotPop_4 : _GEN_3652; // @[Conditional.scala 39:67]
  wire  _GEN_3919 = _T_343 ? spriteVisibleReg_6 : _GEN_3653; // @[Conditional.scala 39:67]
  wire  _GEN_3947 = _T_343 ? planetUp : _GEN_3690; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3962 = _T_343 ? 2'h2 : _GEN_3711; // @[Conditional.scala 39:67]
  wire  _GEN_3995 = _T_343 ? show : _GEN_3744; // @[Conditional.scala 39:67]
  wire  _GEN_4004 = _T_343 ? shipInteract : _GEN_3753; // @[Conditional.scala 39:67]
  wire  _GEN_4067 = _T_343 ? spriteVisibleReg_26 : _GEN_3816; // @[Conditional.scala 39:67]
  wire  _GEN_4070 = _T_343 ? spriteVisibleReg_30 : _GEN_3819; // @[Conditional.scala 39:67]
  wire  _GEN_4073 = _T_343 ? spriteVisibleReg_27 : _GEN_3822; // @[Conditional.scala 39:67]
  wire  _GEN_4076 = _T_343 ? spriteVisibleReg_31 : _GEN_3825; // @[Conditional.scala 39:67]
  wire  _GEN_4079 = _T_343 ? spriteVisibleReg_28 : _GEN_3828; // @[Conditional.scala 39:67]
  wire  _GEN_4082 = _T_343 ? spriteVisibleReg_32 : _GEN_3831; // @[Conditional.scala 39:67]
  wire  _GEN_4085 = _T_343 ? spriteVisibleReg_29 : _GEN_3834; // @[Conditional.scala 39:67]
  wire  _GEN_4088 = _T_343 ? spriteVisibleReg_33 : _GEN_3837; // @[Conditional.scala 39:67]
  wire  _GEN_4091 = _T_343 ? spriteVisibleReg_72 : _GEN_3840; // @[Conditional.scala 39:67]
  wire  _GEN_4092 = _T_343 ? spriteVisibleReg_66 : _GEN_3841; // @[Conditional.scala 39:67]
  wire  _GEN_4093 = _T_343 ? spriteVisibleReg_57 : _GEN_3842; // @[Conditional.scala 39:67]
  wire  _GEN_4094 = _T_343 ? spriteVisibleReg_61 : _GEN_3843; // @[Conditional.scala 39:67]
  wire  _GEN_4095 = _T_343 ? spriteVisibleReg_71 : _GEN_3844; // @[Conditional.scala 39:67]
  wire  _GEN_4096 = _T_343 ? spriteVisibleReg_65 : _GEN_3845; // @[Conditional.scala 39:67]
  wire  _GEN_4097 = _T_343 ? spriteVisibleReg_56 : _GEN_3846; // @[Conditional.scala 39:67]
  wire  _GEN_4098 = _T_343 ? spriteVisibleReg_62 : _GEN_3847; // @[Conditional.scala 39:67]
  wire  _GEN_4099 = _T_343 ? spriteVisibleReg_70 : _GEN_3848; // @[Conditional.scala 39:67]
  wire  _GEN_4100 = _T_343 ? spriteVisibleReg_64 : _GEN_3849; // @[Conditional.scala 39:67]
  wire  _GEN_4101 = _T_343 ? spriteVisibleReg_55 : _GEN_3850; // @[Conditional.scala 39:67]
  wire  _GEN_4102 = _T_343 ? spriteVisibleReg_63 : _GEN_3851; // @[Conditional.scala 39:67]
  wire  _GEN_4103 = _T_343 ? spriteVisibleReg_44 : _GEN_3852; // @[Conditional.scala 39:67]
  wire  _GEN_4106 = _T_343 ? spriteVisibleReg_45 : _GEN_3855; // @[Conditional.scala 39:67]
  wire  _GEN_4109 = _T_343 ? spriteVisibleReg_46 : _GEN_3858; // @[Conditional.scala 39:67]
  wire  _GEN_4112 = _T_343 ? spriteVisibleReg_47 : _GEN_3861; // @[Conditional.scala 39:67]
  wire  _GEN_4115 = _T_343 ? spriteVisibleReg_48 : _GEN_3864; // @[Conditional.scala 39:67]
  wire  _GEN_4118 = _T_343 ? spriteVisibleReg_49 : _GEN_3867; // @[Conditional.scala 39:67]
  wire  _GEN_4121 = _T_343 ? spriteVisibleReg_50 : _GEN_3870; // @[Conditional.scala 39:67]
  wire  _GEN_4124 = _T_343 ? spriteVisibleReg_51 : _GEN_3873; // @[Conditional.scala 39:67]
  wire  _GEN_4127 = _T_343 ? 1'h0 : _GEN_3876; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_4148 = _T_342 ? 6'h0 : _GEN_3897; // @[Conditional.scala 40:58]
  wire [12:0] _GEN_4149 = _T_342 ? 13'h0 : _GEN_3898; // @[Conditional.scala 40:58]
  wire  _GEN_4156 = _T_342 ? shotInteract_0 : _GEN_3905; // @[Conditional.scala 40:58]
  wire  _GEN_4157 = _T_342 ? shotPop_0 : _GEN_3906; // @[Conditional.scala 40:58]
  wire  _GEN_4158 = _T_342 ? spriteVisibleReg_2 : _GEN_3907; // @[Conditional.scala 40:58]
  wire  _GEN_4159 = _T_342 ? shotInteract_1 : _GEN_3908; // @[Conditional.scala 40:58]
  wire  _GEN_4160 = _T_342 ? shotPop_1 : _GEN_3909; // @[Conditional.scala 40:58]
  wire  _GEN_4161 = _T_342 ? spriteVisibleReg_3 : _GEN_3910; // @[Conditional.scala 40:58]
  wire  _GEN_4162 = _T_342 ? shotInteract_2 : _GEN_3911; // @[Conditional.scala 40:58]
  wire  _GEN_4163 = _T_342 ? shotPop_2 : _GEN_3912; // @[Conditional.scala 40:58]
  wire  _GEN_4164 = _T_342 ? spriteVisibleReg_4 : _GEN_3913; // @[Conditional.scala 40:58]
  wire  _GEN_4165 = _T_342 ? shotInteract_3 : _GEN_3914; // @[Conditional.scala 40:58]
  wire  _GEN_4166 = _T_342 ? shotPop_3 : _GEN_3915; // @[Conditional.scala 40:58]
  wire  _GEN_4167 = _T_342 ? spriteVisibleReg_5 : _GEN_3916; // @[Conditional.scala 40:58]
  wire  _GEN_4168 = _T_342 ? shotInteract_4 : _GEN_3917; // @[Conditional.scala 40:58]
  wire  _GEN_4169 = _T_342 ? shotPop_4 : _GEN_3918; // @[Conditional.scala 40:58]
  wire  _GEN_4170 = _T_342 ? spriteVisibleReg_6 : _GEN_3919; // @[Conditional.scala 40:58]
  wire  _GEN_4198 = _T_342 ? planetUp : _GEN_3947; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_4213 = _T_342 ? 2'h2 : _GEN_3962; // @[Conditional.scala 40:58]
  wire  _GEN_4246 = _T_342 ? show : _GEN_3995; // @[Conditional.scala 40:58]
  wire  _GEN_4255 = _T_342 ? shipInteract : _GEN_4004; // @[Conditional.scala 40:58]
  wire  _GEN_4318 = _T_342 ? spriteVisibleReg_26 : _GEN_4067; // @[Conditional.scala 40:58]
  wire  _GEN_4321 = _T_342 ? spriteVisibleReg_30 : _GEN_4070; // @[Conditional.scala 40:58]
  wire  _GEN_4324 = _T_342 ? spriteVisibleReg_27 : _GEN_4073; // @[Conditional.scala 40:58]
  wire  _GEN_4327 = _T_342 ? spriteVisibleReg_31 : _GEN_4076; // @[Conditional.scala 40:58]
  wire  _GEN_4330 = _T_342 ? spriteVisibleReg_28 : _GEN_4079; // @[Conditional.scala 40:58]
  wire  _GEN_4333 = _T_342 ? spriteVisibleReg_32 : _GEN_4082; // @[Conditional.scala 40:58]
  wire  _GEN_4336 = _T_342 ? spriteVisibleReg_29 : _GEN_4085; // @[Conditional.scala 40:58]
  wire  _GEN_4339 = _T_342 ? spriteVisibleReg_33 : _GEN_4088; // @[Conditional.scala 40:58]
  wire  _GEN_4342 = _T_342 ? spriteVisibleReg_72 : _GEN_4091; // @[Conditional.scala 40:58]
  wire  _GEN_4343 = _T_342 ? spriteVisibleReg_66 : _GEN_4092; // @[Conditional.scala 40:58]
  wire  _GEN_4344 = _T_342 ? spriteVisibleReg_57 : _GEN_4093; // @[Conditional.scala 40:58]
  wire  _GEN_4345 = _T_342 ? spriteVisibleReg_61 : _GEN_4094; // @[Conditional.scala 40:58]
  wire  _GEN_4346 = _T_342 ? spriteVisibleReg_71 : _GEN_4095; // @[Conditional.scala 40:58]
  wire  _GEN_4347 = _T_342 ? spriteVisibleReg_65 : _GEN_4096; // @[Conditional.scala 40:58]
  wire  _GEN_4348 = _T_342 ? spriteVisibleReg_56 : _GEN_4097; // @[Conditional.scala 40:58]
  wire  _GEN_4349 = _T_342 ? spriteVisibleReg_62 : _GEN_4098; // @[Conditional.scala 40:58]
  wire  _GEN_4350 = _T_342 ? spriteVisibleReg_70 : _GEN_4099; // @[Conditional.scala 40:58]
  wire  _GEN_4351 = _T_342 ? spriteVisibleReg_64 : _GEN_4100; // @[Conditional.scala 40:58]
  wire  _GEN_4352 = _T_342 ? spriteVisibleReg_55 : _GEN_4101; // @[Conditional.scala 40:58]
  wire  _GEN_4353 = _T_342 ? spriteVisibleReg_63 : _GEN_4102; // @[Conditional.scala 40:58]
  wire  _GEN_4354 = _T_342 ? spriteVisibleReg_44 : _GEN_4103; // @[Conditional.scala 40:58]
  wire  _GEN_4357 = _T_342 ? spriteVisibleReg_45 : _GEN_4106; // @[Conditional.scala 40:58]
  wire  _GEN_4360 = _T_342 ? spriteVisibleReg_46 : _GEN_4109; // @[Conditional.scala 40:58]
  wire  _GEN_4363 = _T_342 ? spriteVisibleReg_47 : _GEN_4112; // @[Conditional.scala 40:58]
  wire  _GEN_4366 = _T_342 ? spriteVisibleReg_48 : _GEN_4115; // @[Conditional.scala 40:58]
  wire  _GEN_4369 = _T_342 ? spriteVisibleReg_49 : _GEN_4118; // @[Conditional.scala 40:58]
  wire  _GEN_4372 = _T_342 ? spriteVisibleReg_50 : _GEN_4121; // @[Conditional.scala 40:58]
  wire  _GEN_4375 = _T_342 ? spriteVisibleReg_51 : _GEN_4124; // @[Conditional.scala 40:58]
  BoxDetection boxDetection ( // @[GameLogic.scala 712:28]
    .clock(boxDetection_clock),
    .io_boxXPosition_0(boxDetection_io_boxXPosition_0),
    .io_boxXPosition_2(boxDetection_io_boxXPosition_2),
    .io_boxXPosition_3(boxDetection_io_boxXPosition_3),
    .io_boxXPosition_4(boxDetection_io_boxXPosition_4),
    .io_boxXPosition_5(boxDetection_io_boxXPosition_5),
    .io_boxXPosition_6(boxDetection_io_boxXPosition_6),
    .io_boxXPosition_7(boxDetection_io_boxXPosition_7),
    .io_boxXPosition_8(boxDetection_io_boxXPosition_8),
    .io_boxXPosition_9(boxDetection_io_boxXPosition_9),
    .io_boxXPosition_10(boxDetection_io_boxXPosition_10),
    .io_boxXPosition_11(boxDetection_io_boxXPosition_11),
    .io_boxXPosition_12(boxDetection_io_boxXPosition_12),
    .io_boxXPosition_13(boxDetection_io_boxXPosition_13),
    .io_boxXPosition_14(boxDetection_io_boxXPosition_14),
    .io_boxXPosition_15(boxDetection_io_boxXPosition_15),
    .io_boxXPosition_16(boxDetection_io_boxXPosition_16),
    .io_boxXPosition_17(boxDetection_io_boxXPosition_17),
    .io_boxYPosition_0(boxDetection_io_boxYPosition_0),
    .io_boxYPosition_2(boxDetection_io_boxYPosition_2),
    .io_boxYPosition_3(boxDetection_io_boxYPosition_3),
    .io_boxYPosition_4(boxDetection_io_boxYPosition_4),
    .io_boxYPosition_5(boxDetection_io_boxYPosition_5),
    .io_boxYPosition_6(boxDetection_io_boxYPosition_6),
    .io_boxYPosition_7(boxDetection_io_boxYPosition_7),
    .io_boxYPosition_8(boxDetection_io_boxYPosition_8),
    .io_boxYPosition_9(boxDetection_io_boxYPosition_9),
    .io_boxYPosition_10(boxDetection_io_boxYPosition_10),
    .io_boxYPosition_11(boxDetection_io_boxYPosition_11),
    .io_boxYPosition_12(boxDetection_io_boxYPosition_12),
    .io_boxYPosition_13(boxDetection_io_boxYPosition_13),
    .io_boxYPosition_14(boxDetection_io_boxYPosition_14),
    .io_boxYPosition_15(boxDetection_io_boxYPosition_15),
    .io_boxYPosition_16(boxDetection_io_boxYPosition_16),
    .io_boxYPosition_17(boxDetection_io_boxYPosition_17),
    .io_overlap_0_7(boxDetection_io_overlap_0_7),
    .io_overlap_0_8(boxDetection_io_overlap_0_8),
    .io_overlap_0_9(boxDetection_io_overlap_0_9),
    .io_overlap_0_10(boxDetection_io_overlap_0_10),
    .io_overlap_0_11(boxDetection_io_overlap_0_11),
    .io_overlap_0_12(boxDetection_io_overlap_0_12),
    .io_overlap_0_13(boxDetection_io_overlap_0_13),
    .io_overlap_0_14(boxDetection_io_overlap_0_14),
    .io_overlap_0_15(boxDetection_io_overlap_0_15),
    .io_overlap_0_16(boxDetection_io_overlap_0_16),
    .io_overlap_0_17(boxDetection_io_overlap_0_17),
    .io_overlap_2_7(boxDetection_io_overlap_2_7),
    .io_overlap_2_8(boxDetection_io_overlap_2_8),
    .io_overlap_2_9(boxDetection_io_overlap_2_9),
    .io_overlap_2_10(boxDetection_io_overlap_2_10),
    .io_overlap_2_11(boxDetection_io_overlap_2_11),
    .io_overlap_2_12(boxDetection_io_overlap_2_12),
    .io_overlap_2_13(boxDetection_io_overlap_2_13),
    .io_overlap_2_14(boxDetection_io_overlap_2_14),
    .io_overlap_2_15(boxDetection_io_overlap_2_15),
    .io_overlap_2_16(boxDetection_io_overlap_2_16),
    .io_overlap_2_17(boxDetection_io_overlap_2_17),
    .io_overlap_3_7(boxDetection_io_overlap_3_7),
    .io_overlap_3_8(boxDetection_io_overlap_3_8),
    .io_overlap_3_9(boxDetection_io_overlap_3_9),
    .io_overlap_3_10(boxDetection_io_overlap_3_10),
    .io_overlap_3_11(boxDetection_io_overlap_3_11),
    .io_overlap_3_12(boxDetection_io_overlap_3_12),
    .io_overlap_3_13(boxDetection_io_overlap_3_13),
    .io_overlap_3_14(boxDetection_io_overlap_3_14),
    .io_overlap_3_15(boxDetection_io_overlap_3_15),
    .io_overlap_3_16(boxDetection_io_overlap_3_16),
    .io_overlap_3_17(boxDetection_io_overlap_3_17),
    .io_overlap_4_7(boxDetection_io_overlap_4_7),
    .io_overlap_4_8(boxDetection_io_overlap_4_8),
    .io_overlap_4_9(boxDetection_io_overlap_4_9),
    .io_overlap_4_10(boxDetection_io_overlap_4_10),
    .io_overlap_4_11(boxDetection_io_overlap_4_11),
    .io_overlap_4_12(boxDetection_io_overlap_4_12),
    .io_overlap_4_13(boxDetection_io_overlap_4_13),
    .io_overlap_4_14(boxDetection_io_overlap_4_14),
    .io_overlap_4_15(boxDetection_io_overlap_4_15),
    .io_overlap_4_16(boxDetection_io_overlap_4_16),
    .io_overlap_4_17(boxDetection_io_overlap_4_17),
    .io_overlap_5_7(boxDetection_io_overlap_5_7),
    .io_overlap_5_8(boxDetection_io_overlap_5_8),
    .io_overlap_5_9(boxDetection_io_overlap_5_9),
    .io_overlap_5_10(boxDetection_io_overlap_5_10),
    .io_overlap_5_11(boxDetection_io_overlap_5_11),
    .io_overlap_5_12(boxDetection_io_overlap_5_12),
    .io_overlap_5_13(boxDetection_io_overlap_5_13),
    .io_overlap_5_14(boxDetection_io_overlap_5_14),
    .io_overlap_5_15(boxDetection_io_overlap_5_15),
    .io_overlap_5_16(boxDetection_io_overlap_5_16),
    .io_overlap_5_17(boxDetection_io_overlap_5_17),
    .io_overlap_6_7(boxDetection_io_overlap_6_7),
    .io_overlap_6_8(boxDetection_io_overlap_6_8),
    .io_overlap_6_9(boxDetection_io_overlap_6_9),
    .io_overlap_6_10(boxDetection_io_overlap_6_10),
    .io_overlap_6_11(boxDetection_io_overlap_6_11),
    .io_overlap_6_12(boxDetection_io_overlap_6_12),
    .io_overlap_6_13(boxDetection_io_overlap_6_13),
    .io_overlap_6_14(boxDetection_io_overlap_6_14),
    .io_overlap_6_15(boxDetection_io_overlap_6_15),
    .io_overlap_6_17(boxDetection_io_overlap_6_17)
  );
  Randomizer Randomizer ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_clock),
    .reset(Randomizer_reset),
    .io_out(Randomizer_io_out)
  );
  Randomizer_1 Randomizer_1 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_1_clock),
    .reset(Randomizer_1_reset),
    .io_out(Randomizer_1_io_out)
  );
  Randomizer_2 Randomizer_2 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_2_clock),
    .reset(Randomizer_2_reset),
    .io_out(Randomizer_2_io_out)
  );
  Randomizer_3 Randomizer_3 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_3_clock),
    .reset(Randomizer_3_reset),
    .io_out(Randomizer_3_io_out)
  );
  Randomizer_4 Randomizer_4 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_4_clock),
    .reset(Randomizer_4_reset),
    .io_out(Randomizer_4_io_out)
  );
  Randomizer_5 Randomizer_5 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_5_clock),
    .reset(Randomizer_5_reset),
    .io_out(Randomizer_5_io_out)
  );
  Randomizer_6 Randomizer_6 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_6_clock),
    .reset(Randomizer_6_reset),
    .io_out(Randomizer_6_io_out)
  );
  Randomizer_7 Randomizer_7 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_7_clock),
    .reset(Randomizer_7_reset),
    .io_out(Randomizer_7_io_out)
  );
  Randomizer_8 Randomizer_8 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_8_clock),
    .reset(Randomizer_8_reset),
    .io_out(Randomizer_8_io_out)
  );
  Randomizer_9 Randomizer_9 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_9_clock),
    .reset(Randomizer_9_reset),
    .io_out(Randomizer_9_io_out)
  );
  Randomizer_10 Randomizer_10 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_10_clock),
    .reset(Randomizer_10_reset),
    .io_out(Randomizer_10_io_out)
  );
  Randomizer_11 Randomizer_11 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_11_clock),
    .reset(Randomizer_11_reset),
    .io_out(Randomizer_11_io_out)
  );
  Randomizer_12 Randomizer_12 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_12_clock),
    .reset(Randomizer_12_reset),
    .io_out(Randomizer_12_io_out)
  );
  Randomizer_13 Randomizer_13 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_13_clock),
    .reset(Randomizer_13_reset),
    .io_out(Randomizer_13_io_out)
  );
  Randomizer_14 Randomizer_14 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_14_clock),
    .reset(Randomizer_14_reset),
    .io_out(Randomizer_14_io_out)
  );
  Randomizer_15 Randomizer_15 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_15_clock),
    .reset(Randomizer_15_reset),
    .io_out(Randomizer_15_io_out)
  );
  Randomizer_16 Randomizer_16 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_16_clock),
    .reset(Randomizer_16_reset),
    .io_out(Randomizer_16_io_out)
  );
  Randomizer_17 Randomizer_17 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_17_clock),
    .reset(Randomizer_17_reset),
    .io_out(Randomizer_17_io_out)
  );
  Randomizer_18 Randomizer_18 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_18_clock),
    .reset(Randomizer_18_reset),
    .io_out(Randomizer_18_io_out)
  );
  Randomizer_19 Randomizer_19 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_19_clock),
    .reset(Randomizer_19_reset),
    .io_out(Randomizer_19_io_out)
  );
  Randomizer Randomizer_20 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_20_clock),
    .reset(Randomizer_20_reset),
    .io_out(Randomizer_20_io_out)
  );
  Randomizer_1 Randomizer_21 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_21_clock),
    .reset(Randomizer_21_reset),
    .io_out(Randomizer_21_io_out)
  );
  Randomizer_2 Randomizer_22 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_22_clock),
    .reset(Randomizer_22_reset),
    .io_out(Randomizer_22_io_out)
  );
  Randomizer_3 Randomizer_23 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_23_clock),
    .reset(Randomizer_23_reset),
    .io_out(Randomizer_23_io_out)
  );
  Randomizer_4 Randomizer_24 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_24_clock),
    .reset(Randomizer_24_reset),
    .io_out(Randomizer_24_io_out)
  );
  Randomizer_5 Randomizer_25 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_25_clock),
    .reset(Randomizer_25_reset),
    .io_out(Randomizer_25_io_out)
  );
  Randomizer_8 Randomizer_26 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_26_clock),
    .reset(Randomizer_26_reset),
    .io_out(Randomizer_26_io_out)
  );
  Randomizer_9 Randomizer_27 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_27_clock),
    .reset(Randomizer_27_reset),
    .io_out(Randomizer_27_io_out)
  );
  Randomizer_10 Randomizer_28 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_28_clock),
    .reset(Randomizer_28_reset),
    .io_out(Randomizer_28_io_out)
  );
  Randomizer_11 Randomizer_29 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_29_clock),
    .reset(Randomizer_29_reset),
    .io_out(Randomizer_29_io_out)
  );
  Randomizer_18 Randomizer_30 ( // @[GameLogic.scala 201:24]
    .clock(Randomizer_30_clock),
    .reset(Randomizer_30_reset),
    .io_out(Randomizer_30_io_out)
  );
  Randomizer_19 Randomizer_31 ( // @[GameLogic.scala 202:31]
    .clock(Randomizer_31_clock),
    .reset(Randomizer_31_reset),
    .io_out(Randomizer_31_io_out)
  );
  Randomizer_4 Randomizer_32 ( // @[GameLogic.scala 374:24]
    .clock(Randomizer_32_clock),
    .reset(Randomizer_32_reset),
    .io_out(Randomizer_32_io_out)
  );
  Randomizer_33 Randomizer_33 ( // @[GameLogic.scala 130:24]
    .clock(Randomizer_33_clock),
    .reset(Randomizer_33_reset),
    .io_out(Randomizer_33_io_out)
  );
  Randomizer_34 Randomizer_34 ( // @[GameLogic.scala 107:24]
    .clock(Randomizer_34_clock),
    .reset(Randomizer_34_reset),
    .io_out(Randomizer_34_io_out)
  );
  Randomizer_35 Randomizer_35 ( // @[GameLogic.scala 108:25]
    .clock(Randomizer_35_clock),
    .reset(Randomizer_35_reset),
    .io_out(Randomizer_35_io_out)
  );
  Randomizer_36 Randomizer_36 ( // @[GameLogic.scala 107:24]
    .clock(Randomizer_36_clock),
    .reset(Randomizer_36_reset),
    .io_out(Randomizer_36_io_out)
  );
  Randomizer_35 Randomizer_37 ( // @[GameLogic.scala 108:25]
    .clock(Randomizer_37_clock),
    .reset(Randomizer_37_reset),
    .io_out(Randomizer_37_io_out)
  );
  Randomizer_38 Randomizer_38 ( // @[GameLogic.scala 107:24]
    .clock(Randomizer_38_clock),
    .reset(Randomizer_38_reset),
    .io_out(Randomizer_38_io_out)
  );
  Randomizer_35 Randomizer_39 ( // @[GameLogic.scala 108:25]
    .clock(Randomizer_39_clock),
    .reset(Randomizer_39_reset),
    .io_out(Randomizer_39_io_out)
  );
  Randomizer_40 Randomizer_40 ( // @[GameLogic.scala 130:24]
    .clock(Randomizer_40_clock),
    .reset(Randomizer_40_reset),
    .io_out(Randomizer_40_io_out)
  );
  Randomizer_41 Randomizer_41 ( // @[GameLogic.scala 107:24]
    .clock(Randomizer_41_clock),
    .reset(Randomizer_41_reset),
    .io_out(Randomizer_41_io_out)
  );
  Randomizer_35 Randomizer_42 ( // @[GameLogic.scala 108:25]
    .clock(Randomizer_42_clock),
    .reset(Randomizer_42_reset),
    .io_out(Randomizer_42_io_out)
  );
  Randomizer_43 Randomizer_43 ( // @[GameLogic.scala 107:24]
    .clock(Randomizer_43_clock),
    .reset(Randomizer_43_reset),
    .io_out(Randomizer_43_io_out)
  );
  Randomizer_35 Randomizer_44 ( // @[GameLogic.scala 108:25]
    .clock(Randomizer_44_clock),
    .reset(Randomizer_44_reset),
    .io_out(Randomizer_44_io_out)
  );
  Randomizer_45 Randomizer_45 ( // @[GameLogic.scala 107:24]
    .clock(Randomizer_45_clock),
    .reset(Randomizer_45_reset),
    .io_out(Randomizer_45_io_out)
  );
  Randomizer_35 Randomizer_46 ( // @[GameLogic.scala 108:25]
    .clock(Randomizer_46_clock),
    .reset(Randomizer_46_reset),
    .io_out(Randomizer_46_io_out)
  );
  assign io_songInput = {{2'd0}, _GEN_4213}; // @[GameLogic.scala 57:16 GameLogic.scala 233:21 GameLogic.scala 233:21 GameLogic.scala 233:21]
  assign io_spriteXPosition_0 = Xstart_0; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_1 = Xstart_1; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_2 = Xstart_2; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_3 = Xstart_3; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_4 = Xstart_4; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_5 = Xstart_5; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_6 = Xstart_6; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_7 = Xstart_7; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_8 = Xstart_8; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_9 = Xstart_9; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_10 = Xstart_10; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_11 = Xstart_11; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_12 = Xstart_12; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_13 = Xstart_13; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_14 = Xstart_14; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_15 = Xstart_15; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_16 = Xstart_16; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_17 = Xstart_17; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_18 = Xstart_18; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_19 = Xstart_19; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_20 = Xstart_20; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_21 = Xstart_21; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_22 = Xstart_22; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_23 = Xstart_23; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_24 = Xstart_24; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_25 = Xstart_25; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_26 = Xstart_26; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_27 = Xstart_27; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_28 = Xstart_28; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_29 = Xstart_29; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_30 = Xstart_30; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_31 = Xstart_31; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_32 = Xstart_32; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_33 = Xstart_33; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_41 = Xstart_41; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_42 = Xstart_42; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_43 = Xstart_43; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_44 = Xstart_44; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_45 = Xstart_45; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_46 = Xstart_46; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_47 = Xstart_47; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_48 = Xstart_48; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_49 = Xstart_49; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_50 = Xstart_50; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_51 = Xstart_51; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_122 = Xstart_122; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_123 = Xstart_123; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_124 = Xstart_124; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_125 = Xstart_125; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_126 = Xstart_126; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteXPosition_127 = Xstart_127; // @[GameLogic.scala 65:21 GameLogic.scala 639:27]
  assign io_spriteYPosition_0 = Ystart_0[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_1 = Ystart_1[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_2 = Ystart_2[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_3 = Ystart_3[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_4 = Ystart_4[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_5 = Ystart_5[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_6 = Ystart_6[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_7 = Ystart_7[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_8 = Ystart_8[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_9 = Ystart_9[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_10 = Ystart_10[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_11 = Ystart_11[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_12 = Ystart_12[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_13 = Ystart_13[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_14 = Ystart_14[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_15 = Ystart_15[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_16 = Ystart_16[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_17 = Ystart_17[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_18 = Ystart_18[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_19 = Ystart_19[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_20 = Ystart_20[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_21 = Ystart_21[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_22 = Ystart_22[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_23 = Ystart_23[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_24 = Ystart_24[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_25 = Ystart_25[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_26 = Ystart_26[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_27 = Ystart_27[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_28 = Ystart_28[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_29 = Ystart_29[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_30 = Ystart_30[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_31 = Ystart_31[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_32 = Ystart_32[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_33 = Ystart_33[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_41 = Ystart_41[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_42 = Ystart_42[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_43 = Ystart_43[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_122 = Ystart_122[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_123 = Ystart_123[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_124 = Ystart_124[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_125 = Ystart_125[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_126 = Ystart_126[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteYPosition_127 = Ystart_127[9:0]; // @[GameLogic.scala 66:22 GameLogic.scala 640:27]
  assign io_spriteVisible_0 = _T_282 ? 1'h0 : spriteVisibleReg_0; // @[GameLogic.scala 67:20 GameLogic.scala 641:25 GameLogic.scala 343:27]
  assign io_spriteVisible_1 = _T_282 ? 1'h0 : spriteVisibleReg_1; // @[GameLogic.scala 67:20 GameLogic.scala 641:25 GameLogic.scala 344:27]
  assign io_spriteVisible_2 = spriteVisibleReg_2; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_3 = spriteVisibleReg_3; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_4 = spriteVisibleReg_4; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_5 = spriteVisibleReg_5; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_6 = spriteVisibleReg_6; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_7 = spriteVisibleReg_7; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_8 = spriteVisibleReg_8; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_9 = spriteVisibleReg_9; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_10 = spriteVisibleReg_10; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_11 = spriteVisibleReg_11; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_12 = spriteVisibleReg_12; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_13 = spriteVisibleReg_13; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_14 = spriteVisibleReg_14; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_15 = spriteVisibleReg_15; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_16 = spriteVisibleReg_16; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_17 = spriteVisibleReg_17; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_18 = spriteVisibleReg_18; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_19 = spriteVisibleReg_19; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_20 = spriteVisibleReg_20; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_21 = spriteVisibleReg_21; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_22 = spriteVisibleReg_22; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_23 = spriteVisibleReg_23; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_24 = spriteVisibleReg_24; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_25 = spriteVisibleReg_25; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_26 = spriteVisibleReg_26; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_27 = spriteVisibleReg_27; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_28 = spriteVisibleReg_28; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_29 = spriteVisibleReg_29; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_30 = spriteVisibleReg_30; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_31 = spriteVisibleReg_31; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_32 = spriteVisibleReg_32; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_33 = spriteVisibleReg_33; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_41 = spriteVisibleReg_41; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_42 = spriteVisibleReg_42; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_43 = spriteVisibleReg_43; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_44 = spriteVisibleReg_44; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_45 = spriteVisibleReg_45; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_46 = spriteVisibleReg_46; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_47 = spriteVisibleReg_47; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_48 = spriteVisibleReg_48; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_49 = spriteVisibleReg_49; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_50 = spriteVisibleReg_50; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_51 = spriteVisibleReg_51; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_55 = spriteVisibleReg_55; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_56 = spriteVisibleReg_56; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_57 = spriteVisibleReg_57; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_61 = spriteVisibleReg_61; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_62 = spriteVisibleReg_62; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_63 = spriteVisibleReg_63; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_64 = spriteVisibleReg_64; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_65 = spriteVisibleReg_65; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_66 = spriteVisibleReg_66; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_70 = spriteVisibleReg_70; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_71 = spriteVisibleReg_71; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteVisible_72 = spriteVisibleReg_72; // @[GameLogic.scala 67:20 GameLogic.scala 641:25]
  assign io_spriteFlipVertical_122 = spriteFlipVerticalReg_122; // @[GameLogic.scala 69:25 GameLogic.scala 643:30]
  assign io_spriteFlipVertical_123 = spriteFlipVerticalReg_123; // @[GameLogic.scala 69:25 GameLogic.scala 643:30]
  assign io_spriteFlipVertical_124 = spriteFlipVerticalReg_124; // @[GameLogic.scala 69:25 GameLogic.scala 643:30]
  assign io_spriteFlipVertical_125 = spriteFlipVerticalReg_125; // @[GameLogic.scala 69:25 GameLogic.scala 643:30]
  assign io_spriteFlipVertical_126 = spriteFlipVerticalReg_126; // @[GameLogic.scala 69:25 GameLogic.scala 643:30]
  assign io_spriteFlipVertical_127 = spriteFlipVerticalReg_127; // @[GameLogic.scala 69:25 GameLogic.scala 643:30]
  assign io_viewBoxX_0 = viewX; // @[GameLogic.scala 645:15 GameLogic.scala 650:18]
  assign io_backBufferWriteData = _GEN_4148[4:0]; // @[GameLogic.scala 654:26 GameLogic.scala 769:36 GameLogic.scala 785:34 GameLogic.scala 799:34 GameLogic.scala 821:34 GameLogic.scala 834:34 GameLogic.scala 848:32]
  assign io_backBufferWriteAddress = _GEN_4149[10:0]; // @[GameLogic.scala 655:29 GameLogic.scala 770:39 GameLogic.scala 786:37 GameLogic.scala 800:37 GameLogic.scala 822:37 GameLogic.scala 835:37 GameLogic.scala 849:35]
  assign io_backBufferWriteEnable = _T_342 ? 1'h0 : _GEN_3899; // @[GameLogic.scala 656:28 GameLogic.scala 771:38 GameLogic.scala 787:36 GameLogic.scala 801:36 GameLogic.scala 823:36 GameLogic.scala 836:36 GameLogic.scala 850:34]
  assign io_frameUpdateDone = _T_342 ? 1'h0 : _GEN_4127; // @[GameLogic.scala 659:22 GameLogic.scala 1037:26]
  assign boxDetection_clock = clock;
  assign boxDetection_io_boxXPosition_0 = $signed(Xstart_0) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_2 = $signed(Xstart_2) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_3 = $signed(Xstart_3) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_4 = $signed(Xstart_4) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_5 = $signed(Xstart_5) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_6 = $signed(Xstart_6) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_7 = $signed(Xstart_7) + $signed(_GEN_4393); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_8 = $signed(Xstart_8) + $signed(_GEN_4395); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_9 = $signed(Xstart_9) + $signed(_GEN_4397); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_10 = $signed(Xstart_10) + $signed(_GEN_4397); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_11 = $signed(Xstart_11) + $signed(_GEN_4397); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_12 = $signed(Xstart_12) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_13 = $signed(Xstart_13) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_14 = $signed(Xstart_14) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_15 = $signed(Xstart_15) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_16 = $signed(Xstart_16) + $signed(_GEN_4379); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxXPosition_17 = $signed(Xstart_17) + $signed(_GEN_4413); // @[GameLogic.scala 714:35]
  assign boxDetection_io_boxYPosition_0 = _T_43[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_2 = _T_71[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_3 = _T_85[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_4 = _T_99[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_5 = _T_113[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_6 = _T_127[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_7 = _T_141[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_8 = _T_155[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_9 = _T_169[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_10 = _T_183[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_11 = _T_197[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_12 = _T_211[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_13 = _T_225[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_14 = _T_239[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_15 = _T_253[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_16 = _T_267[9:0]; // @[GameLogic.scala 715:35]
  assign boxDetection_io_boxYPosition_17 = _T_281[9:0]; // @[GameLogic.scala 715:35]
  assign Randomizer_clock = clock;
  assign Randomizer_reset = reset;
  assign Randomizer_1_clock = clock;
  assign Randomizer_1_reset = reset;
  assign Randomizer_2_clock = clock;
  assign Randomizer_2_reset = reset;
  assign Randomizer_3_clock = clock;
  assign Randomizer_3_reset = reset;
  assign Randomizer_4_clock = clock;
  assign Randomizer_4_reset = reset;
  assign Randomizer_5_clock = clock;
  assign Randomizer_5_reset = reset;
  assign Randomizer_6_clock = clock;
  assign Randomizer_6_reset = reset;
  assign Randomizer_7_clock = clock;
  assign Randomizer_7_reset = reset;
  assign Randomizer_8_clock = clock;
  assign Randomizer_8_reset = reset;
  assign Randomizer_9_clock = clock;
  assign Randomizer_9_reset = reset;
  assign Randomizer_10_clock = clock;
  assign Randomizer_10_reset = reset;
  assign Randomizer_11_clock = clock;
  assign Randomizer_11_reset = reset;
  assign Randomizer_12_clock = clock;
  assign Randomizer_12_reset = reset;
  assign Randomizer_13_clock = clock;
  assign Randomizer_13_reset = reset;
  assign Randomizer_14_clock = clock;
  assign Randomizer_14_reset = reset;
  assign Randomizer_15_clock = clock;
  assign Randomizer_15_reset = reset;
  assign Randomizer_16_clock = clock;
  assign Randomizer_16_reset = reset;
  assign Randomizer_17_clock = clock;
  assign Randomizer_17_reset = reset;
  assign Randomizer_18_clock = clock;
  assign Randomizer_18_reset = reset;
  assign Randomizer_19_clock = clock;
  assign Randomizer_19_reset = reset;
  assign Randomizer_20_clock = clock;
  assign Randomizer_20_reset = reset;
  assign Randomizer_21_clock = clock;
  assign Randomizer_21_reset = reset;
  assign Randomizer_22_clock = clock;
  assign Randomizer_22_reset = reset;
  assign Randomizer_23_clock = clock;
  assign Randomizer_23_reset = reset;
  assign Randomizer_24_clock = clock;
  assign Randomizer_24_reset = reset;
  assign Randomizer_25_clock = clock;
  assign Randomizer_25_reset = reset;
  assign Randomizer_26_clock = clock;
  assign Randomizer_26_reset = reset;
  assign Randomizer_27_clock = clock;
  assign Randomizer_27_reset = reset;
  assign Randomizer_28_clock = clock;
  assign Randomizer_28_reset = reset;
  assign Randomizer_29_clock = clock;
  assign Randomizer_29_reset = reset;
  assign Randomizer_30_clock = clock;
  assign Randomizer_30_reset = reset;
  assign Randomizer_31_clock = clock;
  assign Randomizer_31_reset = reset;
  assign Randomizer_32_clock = clock;
  assign Randomizer_32_reset = reset;
  assign Randomizer_33_clock = clock;
  assign Randomizer_33_reset = reset;
  assign Randomizer_34_clock = clock;
  assign Randomizer_34_reset = reset;
  assign Randomizer_35_clock = clock;
  assign Randomizer_35_reset = reset;
  assign Randomizer_36_clock = clock;
  assign Randomizer_36_reset = reset;
  assign Randomizer_37_clock = clock;
  assign Randomizer_37_reset = reset;
  assign Randomizer_38_clock = clock;
  assign Randomizer_38_reset = reset;
  assign Randomizer_39_clock = clock;
  assign Randomizer_39_reset = reset;
  assign Randomizer_40_clock = clock;
  assign Randomizer_40_reset = reset;
  assign Randomizer_41_clock = clock;
  assign Randomizer_41_reset = reset;
  assign Randomizer_42_clock = clock;
  assign Randomizer_42_reset = reset;
  assign Randomizer_43_clock = clock;
  assign Randomizer_43_reset = reset;
  assign Randomizer_44_clock = clock;
  assign Randomizer_44_reset = reset;
  assign Randomizer_45_clock = clock;
  assign Randomizer_45_reset = reset;
  assign Randomizer_46_clock = clock;
  assign Randomizer_46_reset = reset;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  planetUp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  Xstart_0 = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  Xstart_1 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  Xstart_2 = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  Xstart_3 = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  Xstart_4 = _RAND_5[10:0];
  _RAND_6 = {1{`RANDOM}};
  Xstart_5 = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  Xstart_6 = _RAND_7[10:0];
  _RAND_8 = {1{`RANDOM}};
  Xstart_7 = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  Xstart_8 = _RAND_9[10:0];
  _RAND_10 = {1{`RANDOM}};
  Xstart_9 = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  Xstart_10 = _RAND_11[10:0];
  _RAND_12 = {1{`RANDOM}};
  Xstart_11 = _RAND_12[10:0];
  _RAND_13 = {1{`RANDOM}};
  Xstart_12 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  Xstart_13 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  Xstart_14 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  Xstart_15 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  Xstart_16 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  Xstart_17 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  Xstart_18 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  Xstart_19 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  Xstart_20 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  Xstart_21 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  Xstart_22 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  Xstart_23 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  Xstart_24 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  Xstart_25 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  Xstart_26 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  Xstart_27 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  Xstart_28 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  Xstart_29 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  Xstart_30 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  Xstart_31 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  Xstart_32 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  Xstart_33 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  Xstart_41 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  Xstart_42 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  Xstart_43 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  Xstart_44 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  Xstart_45 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  Xstart_46 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  Xstart_47 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  Xstart_48 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  Xstart_49 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  Xstart_50 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  Xstart_51 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  Xstart_122 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  Xstart_123 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  Xstart_124 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  Xstart_125 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  Xstart_126 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  Xstart_127 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  Ystart_0 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  Ystart_1 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  Ystart_2 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  Ystart_3 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  Ystart_4 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  Ystart_5 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  Ystart_6 = _RAND_58[10:0];
  _RAND_59 = {1{`RANDOM}};
  Ystart_7 = _RAND_59[10:0];
  _RAND_60 = {1{`RANDOM}};
  Ystart_8 = _RAND_60[10:0];
  _RAND_61 = {1{`RANDOM}};
  Ystart_9 = _RAND_61[10:0];
  _RAND_62 = {1{`RANDOM}};
  Ystart_10 = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  Ystart_11 = _RAND_63[10:0];
  _RAND_64 = {1{`RANDOM}};
  Ystart_12 = _RAND_64[10:0];
  _RAND_65 = {1{`RANDOM}};
  Ystart_13 = _RAND_65[10:0];
  _RAND_66 = {1{`RANDOM}};
  Ystart_14 = _RAND_66[10:0];
  _RAND_67 = {1{`RANDOM}};
  Ystart_15 = _RAND_67[10:0];
  _RAND_68 = {1{`RANDOM}};
  Ystart_16 = _RAND_68[10:0];
  _RAND_69 = {1{`RANDOM}};
  Ystart_17 = _RAND_69[10:0];
  _RAND_70 = {1{`RANDOM}};
  Ystart_18 = _RAND_70[10:0];
  _RAND_71 = {1{`RANDOM}};
  Ystart_19 = _RAND_71[10:0];
  _RAND_72 = {1{`RANDOM}};
  Ystart_20 = _RAND_72[10:0];
  _RAND_73 = {1{`RANDOM}};
  Ystart_21 = _RAND_73[10:0];
  _RAND_74 = {1{`RANDOM}};
  Ystart_22 = _RAND_74[10:0];
  _RAND_75 = {1{`RANDOM}};
  Ystart_23 = _RAND_75[10:0];
  _RAND_76 = {1{`RANDOM}};
  Ystart_24 = _RAND_76[10:0];
  _RAND_77 = {1{`RANDOM}};
  Ystart_25 = _RAND_77[10:0];
  _RAND_78 = {1{`RANDOM}};
  Ystart_26 = _RAND_78[10:0];
  _RAND_79 = {1{`RANDOM}};
  Ystart_27 = _RAND_79[10:0];
  _RAND_80 = {1{`RANDOM}};
  Ystart_28 = _RAND_80[10:0];
  _RAND_81 = {1{`RANDOM}};
  Ystart_29 = _RAND_81[10:0];
  _RAND_82 = {1{`RANDOM}};
  Ystart_30 = _RAND_82[10:0];
  _RAND_83 = {1{`RANDOM}};
  Ystart_31 = _RAND_83[10:0];
  _RAND_84 = {1{`RANDOM}};
  Ystart_32 = _RAND_84[10:0];
  _RAND_85 = {1{`RANDOM}};
  Ystart_33 = _RAND_85[10:0];
  _RAND_86 = {1{`RANDOM}};
  Ystart_41 = _RAND_86[10:0];
  _RAND_87 = {1{`RANDOM}};
  Ystart_42 = _RAND_87[10:0];
  _RAND_88 = {1{`RANDOM}};
  Ystart_43 = _RAND_88[10:0];
  _RAND_89 = {1{`RANDOM}};
  Ystart_122 = _RAND_89[10:0];
  _RAND_90 = {1{`RANDOM}};
  Ystart_123 = _RAND_90[10:0];
  _RAND_91 = {1{`RANDOM}};
  Ystart_124 = _RAND_91[10:0];
  _RAND_92 = {1{`RANDOM}};
  Ystart_125 = _RAND_92[10:0];
  _RAND_93 = {1{`RANDOM}};
  Ystart_126 = _RAND_93[10:0];
  _RAND_94 = {1{`RANDOM}};
  Ystart_127 = _RAND_94[10:0];
  _RAND_95 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleReg_32 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleReg_33 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleReg_41 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleReg_42 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleReg_43 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleReg_44 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleReg_45 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleReg_46 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleReg_47 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleReg_48 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleReg_49 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleReg_50 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleReg_51 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleReg_55 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleReg_56 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleReg_57 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleReg_61 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleReg_62 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleReg_63 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleReg_64 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleReg_65 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleReg_66 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleReg_70 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleReg_71 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleReg_72 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteFlipVerticalReg_122 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteFlipVerticalReg_123 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteFlipVerticalReg_124 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteFlipVerticalReg_125 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteFlipVerticalReg_126 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteFlipVerticalReg_127 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  btnCReg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  viewX = _RAND_159[9:0];
  _RAND_160 = {1{`RANDOM}};
  stateReg = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  shotCnt = _RAND_161[9:0];
  _RAND_162 = {1{`RANDOM}};
  shotLoad = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  shotCntBig = _RAND_163[2:0];
  _RAND_164 = {1{`RANDOM}};
  shotCntFast = _RAND_164[2:0];
  _RAND_165 = {1{`RANDOM}};
  shotPop_0 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  shotPop_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  shotPop_2 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  shotPop_3 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  shotPop_4 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  shotInteract_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  shotInteract_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  shotInteract_2 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  shotInteract_3 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  shotInteract_4 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  astInteract_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  astInteract_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  astInteract_2 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  astInteract_3 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  astInteract_4 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  astInteract_5 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  astInteract_6 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  astInteract_7 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  astInteract_8 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  astInteract_9 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  astInteract_10 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  shipInteract = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  die_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  die_1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  die_2 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  die_3 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  die_4 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  die_5 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  die_6 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  die_7 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  die_8 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  die_9 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  die_10 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  kill_0_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  kill_0_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  kill_0_2 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  kill_0_3 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  kill_0_4 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  kill_1_0 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  kill_1_1 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  kill_1_2 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  kill_1_3 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  kill_1_4 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  kill_2_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  kill_2_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  kill_2_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  kill_2_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  kill_2_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  kill_3_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  kill_3_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  kill_3_2 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  kill_3_3 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  kill_3_4 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  kill_4_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  kill_4_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  kill_4_2 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  kill_4_3 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  kill_4_4 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  kill_5_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  kill_5_1 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  kill_5_2 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  kill_5_3 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  kill_5_4 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  kill_6_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  kill_6_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  kill_6_2 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  kill_6_3 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  kill_6_4 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  kill_7_0 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  kill_7_1 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  kill_7_2 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  kill_7_3 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  kill_7_4 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  kill_8_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  kill_8_1 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  kill_8_2 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  kill_8_3 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  kill_8_4 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  kill_9_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  kill_9_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  kill_9_2 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  kill_9_3 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  kill_10_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  kill_10_1 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  kill_10_2 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  kill_10_3 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  kill_10_4 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  hp = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  planetHp = _RAND_253[4:0];
  _RAND_254 = {1{`RANDOM}};
  spwnProt = _RAND_254[5:0];
  _RAND_255 = {1{`RANDOM}};
  show = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  blink = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  secCnt = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  level = _RAND_258[2:0];
  _RAND_259 = {1{`RANDOM}};
  start = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  levelCng = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  cngCnt = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  cnt = _RAND_262[9:0];
  _RAND_263 = {1{`RANDOM}};
  count1 = _RAND_263[6:0];
  _RAND_264 = {1{`RANDOM}};
  count3 = _RAND_264[6:0];
  _RAND_265 = {1{`RANDOM}};
  count4 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  count5 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  _T_913 = _RAND_267[10:0];
  _RAND_268 = {1{`RANDOM}};
  _T_918 = _RAND_268[10:0];
  _RAND_269 = {1{`RANDOM}};
  _T_928 = _RAND_269[10:0];
  _RAND_270 = {1{`RANDOM}};
  _T_933 = _RAND_270[10:0];
  _RAND_271 = {1{`RANDOM}};
  _T_941 = _RAND_271[10:0];
  _RAND_272 = {1{`RANDOM}};
  _T_946 = _RAND_272[10:0];
  _RAND_273 = {1{`RANDOM}};
  _T_954 = _RAND_273[10:0];
  _RAND_274 = {1{`RANDOM}};
  _T_959 = _RAND_274[10:0];
  _RAND_275 = {1{`RANDOM}};
  _T_967 = _RAND_275[10:0];
  _RAND_276 = {1{`RANDOM}};
  _T_972 = _RAND_276[10:0];
  _RAND_277 = {1{`RANDOM}};
  _T_979 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_980 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  _T_981 = _RAND_279[2:0];
  _RAND_280 = {1{`RANDOM}};
  _T_982 = _RAND_280[2:0];
  _RAND_281 = {1{`RANDOM}};
  _T_983 = _RAND_281[2:0];
  _RAND_282 = {1{`RANDOM}};
  _T_1029 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  _T_1030 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_1031 = _RAND_284[2:0];
  _RAND_285 = {1{`RANDOM}};
  _T_1032 = _RAND_285[2:0];
  _RAND_286 = {1{`RANDOM}};
  _T_1033 = _RAND_286[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    planetUp <= reset | _GEN_4198;
    if (reset) begin
      Xstart_0 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (_T_863) begin
                          if (_T_864) begin
                            if (io_btnR) begin
                              if (_T_876) begin
                                Xstart_0 <= _T_879;
                              end
                            end else if (io_btnL) begin
                              if (_T_883) begin
                                Xstart_0 <= _T_886;
                              end
                            end
                          end
                        end else if (!(_T_887)) begin
                          if (_T_978) begin
                            if (die_10) begin
                              if (_T_1135) begin
                                Xstart_0 <= 11'sh40;
                              end else if (die_9) begin
                                if (_T_1135) begin
                                  Xstart_0 <= 11'sh40;
                                end else if (die_8) begin
                                  if (_T_1135) begin
                                    Xstart_0 <= 11'sh40;
                                  end else if (die_7) begin
                                    if (_T_1135) begin
                                      Xstart_0 <= 11'sh40;
                                    end else if (die_6) begin
                                      if (_T_1135) begin
                                        Xstart_0 <= 11'sh40;
                                      end else if (die_5) begin
                                        if (_T_1135) begin
                                          Xstart_0 <= 11'sh40;
                                        end else if (die_4) begin
                                          if (_T_1135) begin
                                            Xstart_0 <= 11'sh40;
                                          end else if (die_3) begin
                                            if (_T_1135) begin
                                              Xstart_0 <= 11'sh40;
                                            end else if (die_2) begin
                                              if (_T_1135) begin
                                                Xstart_0 <= 11'sh40;
                                              end else if (die_1) begin
                                                if (_T_1135) begin
                                                  Xstart_0 <= 11'sh40;
                                                end else if (die_0) begin
                                                  if (_T_1135) begin
                                                    Xstart_0 <= 11'sh40;
                                                  end
                                                end
                                              end else if (die_0) begin
                                                if (_T_1135) begin
                                                  Xstart_0 <= 11'sh40;
                                                end
                                              end
                                            end else if (die_1) begin
                                              if (_T_1135) begin
                                                Xstart_0 <= 11'sh40;
                                              end else if (die_0) begin
                                                if (_T_1135) begin
                                                  Xstart_0 <= 11'sh40;
                                                end
                                              end
                                            end else if (die_0) begin
                                              if (_T_1135) begin
                                                Xstart_0 <= 11'sh40;
                                              end
                                            end
                                          end else if (die_2) begin
                                            if (_T_1135) begin
                                              Xstart_0 <= 11'sh40;
                                            end else if (die_1) begin
                                              if (_T_1135) begin
                                                Xstart_0 <= 11'sh40;
                                              end else begin
                                                Xstart_0 <= _GEN_1182;
                                              end
                                            end else begin
                                              Xstart_0 <= _GEN_1182;
                                            end
                                          end else if (die_1) begin
                                            if (_T_1135) begin
                                              Xstart_0 <= 11'sh40;
                                            end else begin
                                              Xstart_0 <= _GEN_1182;
                                            end
                                          end else begin
                                            Xstart_0 <= _GEN_1182;
                                          end
                                        end else if (die_3) begin
                                          if (_T_1135) begin
                                            Xstart_0 <= 11'sh40;
                                          end else if (die_2) begin
                                            if (_T_1135) begin
                                              Xstart_0 <= 11'sh40;
                                            end else begin
                                              Xstart_0 <= _GEN_1192;
                                            end
                                          end else begin
                                            Xstart_0 <= _GEN_1192;
                                          end
                                        end else if (die_2) begin
                                          if (_T_1135) begin
                                            Xstart_0 <= 11'sh40;
                                          end else begin
                                            Xstart_0 <= _GEN_1192;
                                          end
                                        end else begin
                                          Xstart_0 <= _GEN_1192;
                                        end
                                      end else if (die_4) begin
                                        if (_T_1135) begin
                                          Xstart_0 <= 11'sh40;
                                        end else if (die_3) begin
                                          if (_T_1135) begin
                                            Xstart_0 <= 11'sh40;
                                          end else begin
                                            Xstart_0 <= _GEN_1202;
                                          end
                                        end else begin
                                          Xstart_0 <= _GEN_1202;
                                        end
                                      end else if (die_3) begin
                                        if (_T_1135) begin
                                          Xstart_0 <= 11'sh40;
                                        end else begin
                                          Xstart_0 <= _GEN_1202;
                                        end
                                      end else begin
                                        Xstart_0 <= _GEN_1202;
                                      end
                                    end else if (die_5) begin
                                      if (_T_1135) begin
                                        Xstart_0 <= 11'sh40;
                                      end else if (die_4) begin
                                        if (_T_1135) begin
                                          Xstart_0 <= 11'sh40;
                                        end else begin
                                          Xstart_0 <= _GEN_1212;
                                        end
                                      end else begin
                                        Xstart_0 <= _GEN_1212;
                                      end
                                    end else if (die_4) begin
                                      if (_T_1135) begin
                                        Xstart_0 <= 11'sh40;
                                      end else begin
                                        Xstart_0 <= _GEN_1212;
                                      end
                                    end else begin
                                      Xstart_0 <= _GEN_1212;
                                    end
                                  end else if (die_6) begin
                                    if (_T_1135) begin
                                      Xstart_0 <= 11'sh40;
                                    end else if (die_5) begin
                                      if (_T_1135) begin
                                        Xstart_0 <= 11'sh40;
                                      end else begin
                                        Xstart_0 <= _GEN_1222;
                                      end
                                    end else begin
                                      Xstart_0 <= _GEN_1222;
                                    end
                                  end else if (die_5) begin
                                    if (_T_1135) begin
                                      Xstart_0 <= 11'sh40;
                                    end else begin
                                      Xstart_0 <= _GEN_1222;
                                    end
                                  end else begin
                                    Xstart_0 <= _GEN_1222;
                                  end
                                end else if (die_7) begin
                                  if (_T_1135) begin
                                    Xstart_0 <= 11'sh40;
                                  end else if (die_6) begin
                                    if (_T_1135) begin
                                      Xstart_0 <= 11'sh40;
                                    end else begin
                                      Xstart_0 <= _GEN_1232;
                                    end
                                  end else begin
                                    Xstart_0 <= _GEN_1232;
                                  end
                                end else if (die_6) begin
                                  if (_T_1135) begin
                                    Xstart_0 <= 11'sh40;
                                  end else begin
                                    Xstart_0 <= _GEN_1232;
                                  end
                                end else begin
                                  Xstart_0 <= _GEN_1232;
                                end
                              end else if (die_8) begin
                                if (_T_1135) begin
                                  Xstart_0 <= 11'sh40;
                                end else if (die_7) begin
                                  if (_T_1135) begin
                                    Xstart_0 <= 11'sh40;
                                  end else begin
                                    Xstart_0 <= _GEN_1242;
                                  end
                                end else begin
                                  Xstart_0 <= _GEN_1242;
                                end
                              end else if (die_7) begin
                                if (_T_1135) begin
                                  Xstart_0 <= 11'sh40;
                                end else begin
                                  Xstart_0 <= _GEN_1242;
                                end
                              end else begin
                                Xstart_0 <= _GEN_1242;
                              end
                            end else if (die_9) begin
                              if (_T_1135) begin
                                Xstart_0 <= 11'sh40;
                              end else if (die_8) begin
                                if (_T_1135) begin
                                  Xstart_0 <= 11'sh40;
                                end else begin
                                  Xstart_0 <= _GEN_1252;
                                end
                              end else begin
                                Xstart_0 <= _GEN_1252;
                              end
                            end else if (die_8) begin
                              if (_T_1135) begin
                                Xstart_0 <= 11'sh40;
                              end else begin
                                Xstart_0 <= _GEN_1252;
                              end
                            end else begin
                              Xstart_0 <= _GEN_1252;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_1 <= 11'sh20;
    end else begin
      Xstart_1 <= Xstart_0;
    end
    if (reset) begin
      Xstart_2 <= 11'sh258;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_2 <= _T_349;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (!(_T_706)) begin
                      if (!(_T_863)) begin
                        if (_T_887) begin
                          if (_T_864) begin
                            if (_T_910) begin
                              Xstart_2 <= _T_890;
                            end else if (_T_925) begin
                              Xstart_2 <= _T_890;
                            end else if (shotPop_0) begin
                              if (shotLoad) begin
                                Xstart_2 <= _T_945;
                              end else begin
                                Xstart_2 <= _T_890;
                              end
                            end else begin
                              Xstart_2 <= _T_890;
                            end
                          end else begin
                            Xstart_2 <= _T_890;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_3 <= 11'sh258;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_3 <= _T_352;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (!(_T_706)) begin
                      if (!(_T_863)) begin
                        if (_T_887) begin
                          if (_T_864) begin
                            if (_T_910) begin
                              Xstart_3 <= _T_894;
                            end else if (_T_925) begin
                              Xstart_3 <= _T_894;
                            end else if (shotPop_0) begin
                              Xstart_3 <= _T_894;
                            end else if (shotPop_1) begin
                              if (shotLoad) begin
                                Xstart_3 <= _T_958;
                              end else begin
                                Xstart_3 <= _T_894;
                              end
                            end else begin
                              Xstart_3 <= _T_894;
                            end
                          end else begin
                            Xstart_3 <= _T_894;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_4 <= 11'sh258;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_4 <= _T_355;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (!(_T_706)) begin
                      if (!(_T_863)) begin
                        if (_T_887) begin
                          if (_T_864) begin
                            if (_T_910) begin
                              Xstart_4 <= _T_898;
                            end else if (_T_925) begin
                              Xstart_4 <= _T_898;
                            end else if (shotPop_0) begin
                              Xstart_4 <= _T_898;
                            end else if (shotPop_1) begin
                              Xstart_4 <= _T_898;
                            end else if (shotPop_2) begin
                              if (shotLoad) begin
                                Xstart_4 <= _T_971;
                              end else begin
                                Xstart_4 <= _T_898;
                              end
                            end else begin
                              Xstart_4 <= _T_898;
                            end
                          end else begin
                            Xstart_4 <= _T_898;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_5 <= 11'sh258;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_5 <= _T_358;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (!(_T_706)) begin
                      if (!(_T_863)) begin
                        if (_T_887) begin
                          if (_T_864) begin
                            if (_T_910) begin
                              if (shotPop_3) begin
                                if (shotLoad) begin
                                  Xstart_5 <= _T_917;
                                end else begin
                                  Xstart_5 <= _T_902;
                                end
                              end else begin
                                Xstart_5 <= _T_902;
                              end
                            end else begin
                              Xstart_5 <= _T_902;
                            end
                          end else begin
                            Xstart_5 <= _T_902;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_6 <= 11'sh258;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_6 <= _T_361;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (!(_T_706)) begin
                      if (!(_T_863)) begin
                        if (_T_887) begin
                          if (_T_864) begin
                            if (_T_910) begin
                              Xstart_6 <= _T_906;
                            end else if (_T_925) begin
                              if (shotPop_4) begin
                                if (shotLoad) begin
                                  Xstart_6 <= _T_932;
                                end else begin
                                  Xstart_6 <= _T_906;
                                end
                              end else begin
                                Xstart_6 <= _T_906;
                              end
                            end else begin
                              Xstart_6 <= _T_906;
                            end
                          end else begin
                            Xstart_6 <= _T_906;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_7 <= 11'sh226;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_7 <= _T_364;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (_T_506) begin
              if (_T_508) begin
                if (_T_512) begin
                  if (_T_515) begin
                    if (_T_502) begin
                      Xstart_7 <= _T_295;
                    end else begin
                      Xstart_7 <= _T_526;
                    end
                  end else begin
                    Xstart_7 <= _T_511;
                  end
                end else begin
                  Xstart_7 <= _T_511;
                end
              end
            end else if (!(_T_571)) begin
              if (!(_T_628)) begin
                if (!(_T_685)) begin
                  if (_T_706) begin
                    if (_T_707) begin
                      if (_T_512) begin
                        if (_T_515) begin
                          if (_T_502) begin
                            Xstart_7 <= _T_295;
                          end else begin
                            Xstart_7 <= _T_526;
                          end
                        end else begin
                          Xstart_7 <= _T_511;
                        end
                      end else begin
                        Xstart_7 <= _T_511;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_8 <= 11'sh262;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_8 <= _T_367;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (_T_506) begin
              if (_T_508) begin
                if (_T_512) begin
                  if (_T_533) begin
                    if (_T_502) begin
                      Xstart_8 <= _T_295;
                    end else begin
                      Xstart_8 <= _T_526;
                    end
                  end else begin
                    Xstart_8 <= _T_529;
                  end
                end else begin
                  Xstart_8 <= _T_529;
                end
              end
            end else if (!(_T_571)) begin
              if (!(_T_628)) begin
                if (!(_T_685)) begin
                  if (_T_706) begin
                    if (_T_707) begin
                      if (_T_512) begin
                        if (_T_533) begin
                          if (_T_502) begin
                            Xstart_8 <= _T_295;
                          end else begin
                            Xstart_8 <= _T_526;
                          end
                        end else begin
                          Xstart_8 <= _T_529;
                        end
                      end else begin
                        Xstart_8 <= _T_529;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_9 <= 11'sh320;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_9 <= _T_370;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (_T_506) begin
              if (_T_508) begin
                if (_T_512) begin
                  if (_T_551) begin
                    Xstart_9 <= _GEN_105;
                  end else begin
                    Xstart_9 <= _T_547;
                  end
                end else begin
                  Xstart_9 <= _T_547;
                end
              end
            end else if (!(_T_571)) begin
              if (!(_T_628)) begin
                if (!(_T_685)) begin
                  if (_T_706) begin
                    if (_T_707) begin
                      if (_T_512) begin
                        if (_T_551) begin
                          Xstart_9 <= _GEN_105;
                        end else begin
                          Xstart_9 <= _T_547;
                        end
                      end else begin
                        Xstart_9 <= _T_547;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_10 <= 11'sh320;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_10 <= _T_373;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (_T_571) begin
                if (_T_512) begin
                  if (_T_578) begin
                    Xstart_10 <= _GEN_105;
                  end else begin
                    Xstart_10 <= _T_574;
                  end
                end else begin
                  Xstart_10 <= _T_574;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_11 <= 11'sh2a8;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_11 <= _T_376;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (_T_571) begin
                if (_T_512) begin
                  if (_T_596) begin
                    Xstart_11 <= _GEN_105;
                  end else begin
                    Xstart_11 <= _T_592;
                  end
                end else begin
                  Xstart_11 <= _T_592;
                end
              end else if (!(_T_628)) begin
                if (!(_T_685)) begin
                  if (_T_706) begin
                    if (_T_707) begin
                      if (_T_512) begin
                        if (_T_596) begin
                          Xstart_11 <= _GEN_105;
                        end else begin
                          Xstart_11 <= _T_592;
                        end
                      end else begin
                        Xstart_11 <= _T_592;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_12 <= 11'sh2ee;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_12 <= _T_379;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (_T_571) begin
                if (_T_512) begin
                  if (_T_614) begin
                    Xstart_12 <= _GEN_105;
                  end else begin
                    Xstart_12 <= _T_610;
                  end
                end else begin
                  Xstart_12 <= _T_610;
                end
              end else if (!(_T_628)) begin
                if (!(_T_685)) begin
                  if (_T_706) begin
                    if (_T_707) begin
                      if (_T_512) begin
                        if (_T_614) begin
                          Xstart_12 <= _GEN_105;
                        end else begin
                          Xstart_12 <= _T_610;
                        end
                      end else begin
                        Xstart_12 <= _T_610;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_13 <= 11'sh320;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_13 <= _T_382;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (_T_628) begin
                  if (_T_512) begin
                    if (_T_635) begin
                      Xstart_13 <= _GEN_105;
                    end else begin
                      Xstart_13 <= _T_631;
                    end
                  end else begin
                    Xstart_13 <= _T_631;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_14 <= 11'sh3d4;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_14 <= _T_385;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (_T_628) begin
                  if (_T_512) begin
                    if (_T_653) begin
                      Xstart_14 <= _GEN_105;
                    end else begin
                      Xstart_14 <= _T_649;
                    end
                  end else begin
                    Xstart_14 <= _T_649;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_15 <= 11'sh37a;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_15 <= _T_388;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (_T_628) begin
                  if (_T_512) begin
                    if (_T_671) begin
                      Xstart_15 <= _GEN_105;
                    end else begin
                      Xstart_15 <= _T_667;
                    end
                  end else begin
                    Xstart_15 <= _T_667;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_16 <= 11'sh258;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        Xstart_16 <= _T_391;
      end else if (!(_T_405)) begin
        if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (_T_685) begin
                    if (_T_689) begin
                      if (_T_692) begin
                        Xstart_16 <= _GEN_105;
                      end else begin
                        Xstart_16 <= _T_688;
                      end
                    end else begin
                      Xstart_16 <= _T_688;
                    end
                  end else if (_T_706) begin
                    if (_T_707) begin
                      if (_T_689) begin
                        if (_T_692) begin
                          Xstart_16 <= _GEN_105;
                        end else begin
                          Xstart_16 <= _T_688;
                        end
                      end else begin
                        Xstart_16 <= _T_688;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_17 <= 11'sh80;
    end else if (_T_342) begin
      Xstart_17 <= _T_289;
    end else if (_T_343) begin
      Xstart_17 <= _T_394;
    end else if (_T_405) begin
      Xstart_17 <= _T_289;
    end else if (_T_452) begin
      Xstart_17 <= _T_289;
    end else if (_T_487) begin
      Xstart_17 <= _T_289;
    end else if (_T_506) begin
      Xstart_17 <= _T_289;
    end else if (_T_571) begin
      Xstart_17 <= _T_289;
    end else if (_T_628) begin
      Xstart_17 <= _T_289;
    end else if (_T_685) begin
      Xstart_17 <= _T_289;
    end else if (_T_706) begin
      if (_T_831) begin
        if (_T_834) begin
          Xstart_17 <= _T_526;
        end else if (_T_826) begin
          Xstart_17 <= _T_829;
        end else begin
          Xstart_17 <= 11'sh1e0;
        end
      end else if (_T_826) begin
        Xstart_17 <= _T_829;
      end else begin
        Xstart_17 <= 11'sh1e0;
      end
    end else begin
      Xstart_17 <= _T_289;
    end
    if (reset) begin
      Xstart_18 <= 11'sh60;
    end else begin
      Xstart_18 <= _T_295;
    end
    if (reset) begin
      Xstart_19 <= 11'sh80;
    end else begin
      Xstart_19 <= _T_301;
    end
    if (reset) begin
      Xstart_20 <= 11'sh40;
    end else begin
      Xstart_20 <= _T_289;
    end
    if (reset) begin
      Xstart_21 <= 11'sh60;
    end else begin
      Xstart_21 <= _T_295;
    end
    if (reset) begin
      Xstart_22 <= 11'sh80;
    end else begin
      Xstart_22 <= _T_301;
    end
    if (reset) begin
      Xstart_23 <= 11'sh40;
    end else begin
      Xstart_23 <= _T_289;
    end
    if (reset) begin
      Xstart_24 <= 11'sh60;
    end else begin
      Xstart_24 <= _T_295;
    end
    if (reset) begin
      Xstart_25 <= 11'sh80;
    end else begin
      Xstart_25 <= _T_301;
    end
    if (reset) begin
      Xstart_26 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Xstart_26 <= 11'sh100;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_27 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Xstart_27 <= 11'sh120;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_28 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Xstart_28 <= 11'sh140;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_29 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Xstart_29 <= 11'sh160;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_30 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Xstart_30 <= 11'sh100;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_31 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Xstart_31 <= 11'sh120;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_32 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Xstart_32 <= 11'sh140;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_33 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Xstart_33 <= 11'sh160;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_41 <= 11'sh2bc;
    end else begin
      Xstart_41 <= Xstart_0;
    end
    if (reset) begin
      Xstart_42 <= 11'sh2bc;
    end else begin
      Xstart_42 <= Xstart_0;
    end
    if (reset) begin
      Xstart_43 <= 11'sh2bc;
    end else begin
      Xstart_43 <= Xstart_0;
    end
    if (reset) begin
      Xstart_44 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_44 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_45 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_45 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_46 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_46 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_47 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_47 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_48 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_48 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_49 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_49 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_50 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_50 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_51 <= 11'sh2bc;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              Xstart_51 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_122 <= 11'sh2c0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1043) begin
                                  Xstart_122 <= _T_526;
                                end else begin
                                  Xstart_122 <= _T_1042;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_123 <= 11'sh2c0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1029) begin
                                  if (_T_1058) begin
                                    Xstart_123 <= _T_526;
                                  end else begin
                                    Xstart_123 <= _T_1057;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_124 <= 11'sh2c0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1030) begin
                                  if (_T_1071) begin
                                    Xstart_124 <= _T_526;
                                  end else begin
                                    Xstart_124 <= _T_1070;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_125 <= 11'sh2c0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_993) begin
                                Xstart_125 <= _T_526;
                              end else begin
                                Xstart_125 <= _T_992;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_126 <= 11'sh2c0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_979) begin
                                if (_T_1008) begin
                                  Xstart_126 <= _T_526;
                                end else begin
                                  Xstart_126 <= _T_1007;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_127 <= 11'sh2c0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_980) begin
                                if (_T_1021) begin
                                  Xstart_127 <= _T_526;
                                end else begin
                                  Xstart_127 <= _T_1020;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_0 <= 11'sh148;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (_T_863) begin
                          if (_T_864) begin
                            if (io_btnD) begin
                              if (_T_865) begin
                                Ystart_0 <= _T_868;
                              end
                            end else if (io_btnU) begin
                              if (_T_869) begin
                                Ystart_0 <= _T_872;
                              end
                            end
                          end
                        end else if (!(_T_887)) begin
                          if (_T_978) begin
                            if (die_10) begin
                              if (_T_1135) begin
                                Ystart_0 <= 11'she0;
                              end else if (die_9) begin
                                if (_T_1135) begin
                                  Ystart_0 <= 11'she0;
                                end else if (die_8) begin
                                  if (_T_1135) begin
                                    Ystart_0 <= 11'she0;
                                  end else if (die_7) begin
                                    if (_T_1135) begin
                                      Ystart_0 <= 11'she0;
                                    end else if (die_6) begin
                                      if (_T_1135) begin
                                        Ystart_0 <= 11'she0;
                                      end else if (die_5) begin
                                        if (_T_1135) begin
                                          Ystart_0 <= 11'she0;
                                        end else if (die_4) begin
                                          if (_T_1135) begin
                                            Ystart_0 <= 11'she0;
                                          end else if (die_3) begin
                                            if (_T_1135) begin
                                              Ystart_0 <= 11'she0;
                                            end else if (die_2) begin
                                              if (_T_1135) begin
                                                Ystart_0 <= 11'she0;
                                              end else if (die_1) begin
                                                if (_T_1135) begin
                                                  Ystart_0 <= 11'she0;
                                                end else if (die_0) begin
                                                  if (_T_1135) begin
                                                    Ystart_0 <= 11'she0;
                                                  end
                                                end
                                              end else if (die_0) begin
                                                if (_T_1135) begin
                                                  Ystart_0 <= 11'she0;
                                                end
                                              end
                                            end else if (die_1) begin
                                              if (_T_1135) begin
                                                Ystart_0 <= 11'she0;
                                              end else if (die_0) begin
                                                if (_T_1135) begin
                                                  Ystart_0 <= 11'she0;
                                                end
                                              end
                                            end else if (die_0) begin
                                              if (_T_1135) begin
                                                Ystart_0 <= 11'she0;
                                              end
                                            end
                                          end else if (die_2) begin
                                            if (_T_1135) begin
                                              Ystart_0 <= 11'she0;
                                            end else if (die_1) begin
                                              if (_T_1135) begin
                                                Ystart_0 <= 11'she0;
                                              end else begin
                                                Ystart_0 <= _GEN_1183;
                                              end
                                            end else begin
                                              Ystart_0 <= _GEN_1183;
                                            end
                                          end else if (die_1) begin
                                            if (_T_1135) begin
                                              Ystart_0 <= 11'she0;
                                            end else begin
                                              Ystart_0 <= _GEN_1183;
                                            end
                                          end else begin
                                            Ystart_0 <= _GEN_1183;
                                          end
                                        end else if (die_3) begin
                                          if (_T_1135) begin
                                            Ystart_0 <= 11'she0;
                                          end else if (die_2) begin
                                            if (_T_1135) begin
                                              Ystart_0 <= 11'she0;
                                            end else begin
                                              Ystart_0 <= _GEN_1193;
                                            end
                                          end else begin
                                            Ystart_0 <= _GEN_1193;
                                          end
                                        end else if (die_2) begin
                                          if (_T_1135) begin
                                            Ystart_0 <= 11'she0;
                                          end else begin
                                            Ystart_0 <= _GEN_1193;
                                          end
                                        end else begin
                                          Ystart_0 <= _GEN_1193;
                                        end
                                      end else if (die_4) begin
                                        if (_T_1135) begin
                                          Ystart_0 <= 11'she0;
                                        end else if (die_3) begin
                                          if (_T_1135) begin
                                            Ystart_0 <= 11'she0;
                                          end else begin
                                            Ystart_0 <= _GEN_1203;
                                          end
                                        end else begin
                                          Ystart_0 <= _GEN_1203;
                                        end
                                      end else if (die_3) begin
                                        if (_T_1135) begin
                                          Ystart_0 <= 11'she0;
                                        end else begin
                                          Ystart_0 <= _GEN_1203;
                                        end
                                      end else begin
                                        Ystart_0 <= _GEN_1203;
                                      end
                                    end else if (die_5) begin
                                      if (_T_1135) begin
                                        Ystart_0 <= 11'she0;
                                      end else if (die_4) begin
                                        if (_T_1135) begin
                                          Ystart_0 <= 11'she0;
                                        end else begin
                                          Ystart_0 <= _GEN_1213;
                                        end
                                      end else begin
                                        Ystart_0 <= _GEN_1213;
                                      end
                                    end else if (die_4) begin
                                      if (_T_1135) begin
                                        Ystart_0 <= 11'she0;
                                      end else begin
                                        Ystart_0 <= _GEN_1213;
                                      end
                                    end else begin
                                      Ystart_0 <= _GEN_1213;
                                    end
                                  end else if (die_6) begin
                                    if (_T_1135) begin
                                      Ystart_0 <= 11'she0;
                                    end else if (die_5) begin
                                      if (_T_1135) begin
                                        Ystart_0 <= 11'she0;
                                      end else begin
                                        Ystart_0 <= _GEN_1223;
                                      end
                                    end else begin
                                      Ystart_0 <= _GEN_1223;
                                    end
                                  end else if (die_5) begin
                                    if (_T_1135) begin
                                      Ystart_0 <= 11'she0;
                                    end else begin
                                      Ystart_0 <= _GEN_1223;
                                    end
                                  end else begin
                                    Ystart_0 <= _GEN_1223;
                                  end
                                end else if (die_7) begin
                                  if (_T_1135) begin
                                    Ystart_0 <= 11'she0;
                                  end else if (die_6) begin
                                    if (_T_1135) begin
                                      Ystart_0 <= 11'she0;
                                    end else begin
                                      Ystart_0 <= _GEN_1233;
                                    end
                                  end else begin
                                    Ystart_0 <= _GEN_1233;
                                  end
                                end else if (die_6) begin
                                  if (_T_1135) begin
                                    Ystart_0 <= 11'she0;
                                  end else begin
                                    Ystart_0 <= _GEN_1233;
                                  end
                                end else begin
                                  Ystart_0 <= _GEN_1233;
                                end
                              end else if (die_8) begin
                                if (_T_1135) begin
                                  Ystart_0 <= 11'she0;
                                end else if (die_7) begin
                                  if (_T_1135) begin
                                    Ystart_0 <= 11'she0;
                                  end else begin
                                    Ystart_0 <= _GEN_1243;
                                  end
                                end else begin
                                  Ystart_0 <= _GEN_1243;
                                end
                              end else if (die_7) begin
                                if (_T_1135) begin
                                  Ystart_0 <= 11'she0;
                                end else begin
                                  Ystart_0 <= _GEN_1243;
                                end
                              end else begin
                                Ystart_0 <= _GEN_1243;
                              end
                            end else if (die_9) begin
                              if (_T_1135) begin
                                Ystart_0 <= 11'she0;
                              end else if (die_8) begin
                                if (_T_1135) begin
                                  Ystart_0 <= 11'she0;
                                end else begin
                                  Ystart_0 <= _GEN_1253;
                                end
                              end else begin
                                Ystart_0 <= _GEN_1253;
                              end
                            end else if (die_8) begin
                              if (_T_1135) begin
                                Ystart_0 <= 11'she0;
                              end else begin
                                Ystart_0 <= _GEN_1253;
                              end
                            end else begin
                              Ystart_0 <= _GEN_1253;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_1 <= 11'sh148;
    end else begin
      Ystart_1 <= Ystart_0;
    end
    if (reset) begin
      Ystart_2 <= 11'sh64;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (!(_T_910)) begin
                                if (!(_T_925)) begin
                                  if (shotPop_0) begin
                                    if (shotLoad) begin
                                      Ystart_2 <= _T_946;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_3 <= 11'sh96;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (!(_T_910)) begin
                                if (!(_T_925)) begin
                                  if (!(shotPop_0)) begin
                                    if (shotPop_1) begin
                                      if (shotLoad) begin
                                        Ystart_3 <= _T_959;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_4 <= 11'sh64;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (!(_T_910)) begin
                                if (!(_T_925)) begin
                                  if (!(shotPop_0)) begin
                                    if (!(shotPop_1)) begin
                                      if (shotPop_2) begin
                                        if (shotLoad) begin
                                          Ystart_4 <= _T_972;
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_5 <= 11'sh64;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (_T_910) begin
                                if (shotPop_3) begin
                                  if (shotLoad) begin
                                    Ystart_5 <= _T_918;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_6 <= 11'sh64;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (!(_T_910)) begin
                                if (_T_925) begin
                                  if (shotPop_4) begin
                                    if (shotLoad) begin
                                      Ystart_6 <= _T_933;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_7 <= 11'sh64;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (_T_506) begin
                if (_T_508) begin
                  if (_T_512) begin
                    if (_T_515) begin
                      if (_T_502) begin
                        Ystart_7 <= _T_522;
                      end else begin
                        Ystart_7 <= {{1{Randomizer_io_out[9]}},Randomizer_io_out};
                      end
                    end
                  end
                end
              end else if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (_T_706) begin
                      if (_T_707) begin
                        if (_T_512) begin
                          if (_T_515) begin
                            if (_T_502) begin
                              Ystart_7 <= _T_721;
                            end else begin
                              Ystart_7 <= {{1{Randomizer_20_io_out[9]}},Randomizer_20_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_8 <= 11'sh7d;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (_T_506) begin
                if (_T_508) begin
                  if (_T_512) begin
                    if (_T_533) begin
                      if (_T_502) begin
                        Ystart_8 <= _T_540;
                      end else begin
                        Ystart_8 <= {{1{Randomizer_2_io_out[9]}},Randomizer_2_io_out};
                      end
                    end
                  end
                end
              end else if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (_T_706) begin
                      if (_T_707) begin
                        if (_T_512) begin
                          if (_T_533) begin
                            if (_T_502) begin
                              Ystart_8 <= _T_739;
                            end else begin
                              Ystart_8 <= {{1{Randomizer_22_io_out[9]}},Randomizer_22_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_9 <= 11'sh96;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (_T_506) begin
                if (_T_508) begin
                  if (_T_512) begin
                    if (_T_551) begin
                      if (_T_502) begin
                        Ystart_9 <= _T_558;
                      end else begin
                        Ystart_9 <= {{1{Randomizer_4_io_out[9]}},Randomizer_4_io_out};
                      end
                    end
                  end
                end
              end else if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (_T_706) begin
                      if (_T_707) begin
                        if (_T_512) begin
                          if (_T_551) begin
                            if (_T_502) begin
                              Ystart_9 <= _T_757;
                            end else begin
                              Ystart_9 <= {{1{Randomizer_24_io_out[9]}},Randomizer_24_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_10 <= 11'shaa;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (_T_571) begin
                  if (_T_512) begin
                    if (_T_578) begin
                      if (_T_502) begin
                        Ystart_10 <= _T_585;
                      end else begin
                        Ystart_10 <= {{1{Randomizer_6_io_out[9]}},Randomizer_6_io_out};
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_11 <= 11'shb4;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (_T_571) begin
                  if (_T_512) begin
                    if (_T_596) begin
                      if (_T_502) begin
                        Ystart_11 <= _T_603;
                      end else begin
                        Ystart_11 <= {{1{Randomizer_8_io_out[9]}},Randomizer_8_io_out};
                      end
                    end
                  end
                end else if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (_T_706) begin
                      if (_T_707) begin
                        if (_T_512) begin
                          if (_T_596) begin
                            if (_T_502) begin
                              Ystart_11 <= _T_775;
                            end else begin
                              Ystart_11 <= {{1{Randomizer_26_io_out[9]}},Randomizer_26_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_12 <= 11'shc8;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (_T_571) begin
                  if (_T_512) begin
                    if (_T_614) begin
                      if (_T_502) begin
                        Ystart_12 <= _T_621;
                      end else begin
                        Ystart_12 <= {{1{Randomizer_10_io_out[9]}},Randomizer_10_io_out};
                      end
                    end
                  end
                end else if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (_T_706) begin
                      if (_T_707) begin
                        if (_T_512) begin
                          if (_T_614) begin
                            if (_T_502) begin
                              Ystart_12 <= _T_793;
                            end else begin
                              Ystart_12 <= {{1{Randomizer_28_io_out[9]}},Randomizer_28_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_13 <= 11'shfa;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (_T_628) begin
                    if (_T_512) begin
                      if (_T_635) begin
                        if (_T_502) begin
                          Ystart_13 <= _T_642;
                        end else begin
                          Ystart_13 <= {{1{Randomizer_12_io_out[9]}},Randomizer_12_io_out};
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_14 <= 11'sh12c;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (_T_628) begin
                    if (_T_512) begin
                      if (_T_653) begin
                        if (_T_502) begin
                          Ystart_14 <= _T_660;
                        end else begin
                          Ystart_14 <= {{1{Randomizer_14_io_out[9]}},Randomizer_14_io_out};
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_15 <= 11'sh14c;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (_T_628) begin
                    if (_T_512) begin
                      if (_T_671) begin
                        if (_T_502) begin
                          Ystart_15 <= _T_678;
                        end else begin
                          Ystart_15 <= {{1{Randomizer_16_io_out[9]}},Randomizer_16_io_out};
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_16 <= 11'shc8;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (_T_685) begin
                      if (_T_689) begin
                        if (_T_692) begin
                          if (_T_502) begin
                            Ystart_16 <= _T_699;
                          end else begin
                            Ystart_16 <= {{1{Randomizer_18_io_out[9]}},Randomizer_18_io_out};
                          end
                        end
                      end
                    end else if (_T_706) begin
                      if (_T_707) begin
                        if (_T_689) begin
                          if (_T_692) begin
                            if (_T_502) begin
                              Ystart_16 <= _T_811;
                            end else begin
                              Ystart_16 <= {{1{Randomizer_30_io_out[9]}},Randomizer_30_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_17 <= 11'sh80;
    end else if (_T_342) begin
      Ystart_17 <= _T_292;
    end else if (_T_343) begin
      Ystart_17 <= _T_292;
    end else if (_T_405) begin
      Ystart_17 <= _T_292;
    end else if (_T_452) begin
      Ystart_17 <= _T_292;
    end else if (_T_487) begin
      Ystart_17 <= _T_292;
    end else if (_T_506) begin
      Ystart_17 <= _T_292;
    end else if (_T_571) begin
      Ystart_17 <= _T_292;
    end else if (_T_628) begin
      Ystart_17 <= _T_292;
    end else if (_T_685) begin
      Ystart_17 <= _T_292;
    end else if (_T_706) begin
      if (_T_831) begin
        if (_T_834) begin
          Ystart_17 <= {{1{_T_846[9]}},_T_846};
        end else begin
          Ystart_17 <= _T_825;
        end
      end else begin
        Ystart_17 <= _T_825;
      end
    end else begin
      Ystart_17 <= _T_292;
    end
    if (reset) begin
      Ystart_18 <= 11'sh40;
    end else begin
      Ystart_18 <= _T_292;
    end
    if (reset) begin
      Ystart_19 <= 11'sh40;
    end else begin
      Ystart_19 <= _T_292;
    end
    if (reset) begin
      Ystart_20 <= 11'sh60;
    end else begin
      Ystart_20 <= _T_310;
    end
    if (reset) begin
      Ystart_21 <= 11'sh60;
    end else begin
      Ystart_21 <= _T_310;
    end
    if (reset) begin
      Ystart_22 <= 11'sh60;
    end else begin
      Ystart_22 <= _T_310;
    end
    if (reset) begin
      Ystart_23 <= 11'sh80;
    end else begin
      Ystart_23 <= _T_328;
    end
    if (reset) begin
      Ystart_24 <= 11'sh80;
    end else begin
      Ystart_24 <= _T_328;
    end
    if (reset) begin
      Ystart_25 <= 11'sh80;
    end else begin
      Ystart_25 <= _T_328;
    end
    if (reset) begin
      Ystart_26 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Ystart_26 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_27 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Ystart_27 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_28 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Ystart_28 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_29 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_282) begin
                                Ystart_29 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_30 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Ystart_30 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_31 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Ystart_31 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_32 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Ystart_32 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_33 <= 11'sh20;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_501) begin
                                Ystart_33 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_41 <= 11'sh20;
    end else begin
      Ystart_41 <= Ystart_0;
    end
    if (reset) begin
      Ystart_42 <= 11'sh20;
    end else begin
      Ystart_42 <= Ystart_0;
    end
    if (reset) begin
      Ystart_43 <= 11'sh20;
    end else begin
      Ystart_43 <= Ystart_0;
    end
    if (reset) begin
      Ystart_122 <= 11'sh96;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1043) begin
                                  Ystart_122 <= {{1{Randomizer_41_io_out[9]}},Randomizer_41_io_out};
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_123 <= 11'shfa;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1029) begin
                                  if (_T_1058) begin
                                    Ystart_123 <= {{1{Randomizer_43_io_out[9]}},Randomizer_43_io_out};
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_124 <= 11'sh140;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1030) begin
                                  if (_T_1071) begin
                                    Ystart_124 <= {{1{Randomizer_45_io_out[9]}},Randomizer_45_io_out};
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_125 <= 11'shd2;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_993) begin
                                Ystart_125 <= {{1{Randomizer_34_io_out[9]}},Randomizer_34_io_out};
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_126 <= 11'sh64;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_979) begin
                                if (_T_1008) begin
                                  Ystart_126 <= {{1{Randomizer_36_io_out[9]}},Randomizer_36_io_out};
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_127 <= 11'sh12c;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_980) begin
                                if (_T_1021) begin
                                  Ystart_127 <= {{1{Randomizer_38_io_out[9]}},Randomizer_38_io_out};
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    spriteVisibleReg_0 <= reset | _GEN_0;
    spriteVisibleReg_1 <= reset | _GEN_1;
    spriteVisibleReg_2 <= reset | _GEN_4158;
    spriteVisibleReg_3 <= reset | _GEN_4161;
    spriteVisibleReg_4 <= reset | _GEN_4164;
    spriteVisibleReg_5 <= reset | _GEN_4167;
    spriteVisibleReg_6 <= reset | _GEN_4170;
    if (reset) begin
      spriteVisibleReg_7 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_506) begin
      if (_T_508) begin
        if (kill_0_4) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_3) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_2) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_1) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_0) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_7 <= _GEN_108;
        end else begin
          spriteVisibleReg_7 <= _GEN_9;
        end
      end else begin
        spriteVisibleReg_7 <= _GEN_9;
      end
    end else if (_T_571) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_628) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_685) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_0_4) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_3) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_2) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_1) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_0) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_7 <= _GEN_108;
        end else begin
          spriteVisibleReg_7 <= _GEN_9;
        end
      end else begin
        spriteVisibleReg_7 <= _GEN_9;
      end
    end else if (_T_863) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_887) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_7 <= 1'h0;
      end else begin
        spriteVisibleReg_7 <= _GEN_9;
      end
    end else begin
      spriteVisibleReg_7 <= _GEN_9;
    end
    if (reset) begin
      spriteVisibleReg_8 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_506) begin
      if (_T_508) begin
        if (kill_1_4) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_3) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_2) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_1) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_0) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_8 <= _GEN_158;
        end else begin
          spriteVisibleReg_8 <= _GEN_11;
        end
      end else begin
        spriteVisibleReg_8 <= _GEN_11;
      end
    end else if (_T_571) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_628) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_685) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_1_4) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_3) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_2) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_1) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_0) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_8 <= _GEN_158;
        end else begin
          spriteVisibleReg_8 <= _GEN_11;
        end
      end else begin
        spriteVisibleReg_8 <= _GEN_11;
      end
    end else if (_T_863) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_887) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_8 <= 1'h0;
      end else begin
        spriteVisibleReg_8 <= _GEN_11;
      end
    end else begin
      spriteVisibleReg_8 <= _GEN_11;
    end
    if (reset) begin
      spriteVisibleReg_9 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_506) begin
      if (_T_508) begin
        if (kill_2_4) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_3) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_2) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_1) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_0) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_9 <= _GEN_208;
        end else begin
          spriteVisibleReg_9 <= _GEN_13;
        end
      end else begin
        spriteVisibleReg_9 <= _GEN_13;
      end
    end else if (_T_571) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_628) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_685) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_2_4) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_3) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_2) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_1) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_0) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_9 <= _GEN_208;
        end else begin
          spriteVisibleReg_9 <= _GEN_13;
        end
      end else begin
        spriteVisibleReg_9 <= _GEN_13;
      end
    end else if (_T_863) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_887) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_9 <= 1'h0;
      end else begin
        spriteVisibleReg_9 <= _GEN_13;
      end
    end else begin
      spriteVisibleReg_9 <= _GEN_13;
    end
    if (reset) begin
      spriteVisibleReg_10 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_506) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_571) begin
      if (kill_3_4) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_3) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_2) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_1) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_0) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (_T_512) begin
        spriteVisibleReg_10 <= _GEN_286;
      end else begin
        spriteVisibleReg_10 <= _GEN_15;
      end
    end else if (_T_628) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_685) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_706) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_863) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_887) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_10 <= 1'h0;
      end else begin
        spriteVisibleReg_10 <= _GEN_15;
      end
    end else begin
      spriteVisibleReg_10 <= _GEN_15;
    end
    if (reset) begin
      spriteVisibleReg_11 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_506) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_571) begin
      if (kill_4_4) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_3) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_2) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_1) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_0) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (_T_512) begin
        spriteVisibleReg_11 <= _GEN_336;
      end else begin
        spriteVisibleReg_11 <= _GEN_17;
      end
    end else if (_T_628) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_685) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_4_4) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_3) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_2) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_1) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_0) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_11 <= _GEN_336;
        end else begin
          spriteVisibleReg_11 <= _GEN_17;
        end
      end else begin
        spriteVisibleReg_11 <= _GEN_17;
      end
    end else if (_T_863) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_887) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_11 <= 1'h0;
      end else begin
        spriteVisibleReg_11 <= _GEN_17;
      end
    end else begin
      spriteVisibleReg_11 <= _GEN_17;
    end
    if (reset) begin
      spriteVisibleReg_12 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_506) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_571) begin
      if (kill_5_4) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_3) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_2) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_1) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_0) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (_T_512) begin
        spriteVisibleReg_12 <= _GEN_386;
      end else begin
        spriteVisibleReg_12 <= _GEN_19;
      end
    end else if (_T_628) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_685) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_5_4) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_3) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_2) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_1) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_0) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (_T_512) begin
          spriteVisibleReg_12 <= _GEN_386;
        end else begin
          spriteVisibleReg_12 <= _GEN_19;
        end
      end else begin
        spriteVisibleReg_12 <= _GEN_19;
      end
    end else if (_T_863) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_887) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_12 <= 1'h0;
      end else begin
        spriteVisibleReg_12 <= _GEN_19;
      end
    end else begin
      spriteVisibleReg_12 <= _GEN_19;
    end
    if (reset) begin
      spriteVisibleReg_13 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_506) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_571) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_628) begin
      if (kill_6_4) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_3) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_2) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_1) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_0) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (_T_512) begin
        spriteVisibleReg_13 <= _GEN_436;
      end else begin
        spriteVisibleReg_13 <= _GEN_21;
      end
    end else if (_T_685) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_706) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_863) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_887) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_13 <= 1'h0;
      end else begin
        spriteVisibleReg_13 <= _GEN_21;
      end
    end else begin
      spriteVisibleReg_13 <= _GEN_21;
    end
    if (reset) begin
      spriteVisibleReg_14 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_506) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_571) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_628) begin
      if (kill_7_4) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_3) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_2) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_1) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_0) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (_T_512) begin
        spriteVisibleReg_14 <= _GEN_486;
      end else begin
        spriteVisibleReg_14 <= _GEN_23;
      end
    end else if (_T_685) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_706) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_863) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_887) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_14 <= 1'h0;
      end else begin
        spriteVisibleReg_14 <= _GEN_23;
      end
    end else begin
      spriteVisibleReg_14 <= _GEN_23;
    end
    if (reset) begin
      spriteVisibleReg_15 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_506) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_571) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_628) begin
      if (kill_8_4) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_3) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_2) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_1) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_0) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (_T_512) begin
        spriteVisibleReg_15 <= _GEN_536;
      end else begin
        spriteVisibleReg_15 <= _GEN_25;
      end
    end else if (_T_685) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_706) begin
      spriteVisibleReg_15 <= 1'h0;
    end else if (_T_863) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_887) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_15 <= 1'h0;
      end else begin
        spriteVisibleReg_15 <= _GEN_25;
      end
    end else begin
      spriteVisibleReg_15 <= _GEN_25;
    end
    if (reset) begin
      spriteVisibleReg_16 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_506) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_571) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_628) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_685) begin
      if (kill_9_3) begin
        spriteVisibleReg_16 <= 1'h0;
      end else if (_T_689) begin
        spriteVisibleReg_16 <= _GEN_586;
      end else begin
        spriteVisibleReg_16 <= _GEN_27;
      end
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_9_3) begin
          spriteVisibleReg_16 <= 1'h0;
        end else if (_T_689) begin
          spriteVisibleReg_16 <= _GEN_586;
        end else begin
          spriteVisibleReg_16 <= _GEN_27;
        end
      end else begin
        spriteVisibleReg_16 <= _GEN_27;
      end
    end else if (_T_863) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_887) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_978) begin
      if (_T_1086) begin
        spriteVisibleReg_16 <= 1'h0;
      end else begin
        spriteVisibleReg_16 <= _GEN_27;
      end
    end else begin
      spriteVisibleReg_16 <= _GEN_27;
    end
    if (reset) begin
      spriteVisibleReg_17 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_487) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_506) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_571) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_628) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_685) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_706) begin
      if (_T_501) begin
        spriteVisibleReg_17 <= 1'h0;
      end else if (_T_831) begin
        spriteVisibleReg_17 <= _GEN_827;
      end else begin
        spriteVisibleReg_17 <= _GEN_29;
      end
    end else begin
      spriteVisibleReg_17 <= _GEN_29;
    end
    spriteVisibleReg_18 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_19 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_20 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_21 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_22 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_23 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_24 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_25 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_26 <= reset | _GEN_4318;
    spriteVisibleReg_27 <= reset | _GEN_4324;
    spriteVisibleReg_28 <= reset | _GEN_4330;
    spriteVisibleReg_29 <= reset | _GEN_4336;
    spriteVisibleReg_30 <= reset | _GEN_4321;
    spriteVisibleReg_31 <= reset | _GEN_4327;
    spriteVisibleReg_32 <= reset | _GEN_4333;
    spriteVisibleReg_33 <= reset | _GEN_4339;
    spriteVisibleReg_41 <= reset | _GEN_4;
    spriteVisibleReg_42 <= reset | _GEN_5;
    spriteVisibleReg_43 <= reset | _GEN_6;
    spriteVisibleReg_44 <= reset | _GEN_4354;
    spriteVisibleReg_45 <= reset | _GEN_4357;
    spriteVisibleReg_46 <= reset | _GEN_4360;
    spriteVisibleReg_47 <= reset | _GEN_4363;
    spriteVisibleReg_48 <= reset | _GEN_4366;
    spriteVisibleReg_49 <= reset | _GEN_4369;
    spriteVisibleReg_50 <= reset | _GEN_4372;
    spriteVisibleReg_51 <= reset | _GEN_4375;
    spriteVisibleReg_55 <= reset | _GEN_4352;
    spriteVisibleReg_56 <= reset | _GEN_4348;
    spriteVisibleReg_57 <= reset | _GEN_4344;
    spriteVisibleReg_61 <= reset | _GEN_4345;
    spriteVisibleReg_62 <= reset | _GEN_4349;
    spriteVisibleReg_63 <= reset | _GEN_4353;
    spriteVisibleReg_64 <= reset | _GEN_4351;
    spriteVisibleReg_65 <= reset | _GEN_4347;
    spriteVisibleReg_66 <= reset | _GEN_4343;
    spriteVisibleReg_70 <= reset | _GEN_4350;
    spriteVisibleReg_71 <= reset | _GEN_4346;
    spriteVisibleReg_72 <= reset | _GEN_4342;
    if (reset) begin
      spriteFlipVerticalReg_122 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1043) begin
                                  spriteFlipVerticalReg_122 <= _T_1048;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_123 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1029) begin
                                  if (_T_1058) begin
                                    spriteFlipVerticalReg_123 <= _T_1063;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_124 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1028) begin
                                if (_T_1030) begin
                                  if (_T_1071) begin
                                    spriteFlipVerticalReg_124 <= _T_1076;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_125 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_993) begin
                                spriteFlipVerticalReg_125 <= _T_998;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_126 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_979) begin
                                if (_T_1008) begin
                                  spriteFlipVerticalReg_126 <= _T_1013;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_127 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_980) begin
                                if (_T_1021) begin
                                  spriteFlipVerticalReg_127 <= _T_1026;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btnCReg <= io_btnC;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              btnCReg <= io_btnC;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      viewX <= 10'h0;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        if (_T_396) begin
          viewX <= _T_402;
        end else begin
          viewX <= _T_346;
        end
      end
    end
    if (reset) begin
      stateReg <= 4'h0;
    end else if (_T_342) begin
      if (io_newFrame) begin
        stateReg <= 4'h1;
      end
    end else if (_T_343) begin
      if (levelCng) begin
        stateReg <= 4'h2;
      end else begin
        stateReg <= 4'h5;
      end
    end else if (_T_405) begin
      if (_T_438) begin
        if (_T_409) begin
          stateReg <= 4'h2;
        end else if (_T_424) begin
          if (_T_409) begin
            stateReg <= 4'h2;
          end else if (_T_407) begin
            if (_T_408) begin
              if (_T_409) begin
                stateReg <= 4'h2;
              end else begin
                stateReg <= 4'h3;
              end
            end else begin
              stateReg <= 4'h3;
            end
          end else begin
            stateReg <= 4'h3;
          end
        end else if (_T_407) begin
          if (_T_408) begin
            if (_T_409) begin
              stateReg <= 4'h2;
            end else begin
              stateReg <= 4'h3;
            end
          end else begin
            stateReg <= 4'h3;
          end
        end else begin
          stateReg <= 4'h3;
        end
      end else if (_T_424) begin
        if (_T_409) begin
          stateReg <= 4'h2;
        end else if (_T_407) begin
          if (_T_408) begin
            if (_T_409) begin
              stateReg <= 4'h2;
            end else begin
              stateReg <= 4'h3;
            end
          end else begin
            stateReg <= 4'h3;
          end
        end else begin
          stateReg <= 4'h3;
        end
      end else if (_T_407) begin
        if (_T_408) begin
          if (_T_409) begin
            stateReg <= 4'h2;
          end else begin
            stateReg <= 4'h3;
          end
        end else begin
          stateReg <= 4'h3;
        end
      end else begin
        stateReg <= 4'h3;
      end
    end else if (_T_452) begin
      if (_T_438) begin
        if (_T_409) begin
          stateReg <= 4'h3;
        end else if (_T_424) begin
          if (_T_409) begin
            stateReg <= 4'h3;
          end else begin
            stateReg <= 4'h4;
          end
        end else begin
          stateReg <= 4'h4;
        end
      end else if (_T_424) begin
        if (_T_409) begin
          stateReg <= 4'h3;
        end else begin
          stateReg <= 4'h4;
        end
      end else begin
        stateReg <= 4'h4;
      end
    end else if (_T_487) begin
      if (_T_409) begin
        stateReg <= 4'h4;
      end else if (_T_501) begin
        stateReg <= 4'ha;
      end else if (_T_504) begin
        stateReg <= 4'h9;
      end else begin
        stateReg <= 4'h5;
      end
    end else if (_T_506) begin
      if (_T_508) begin
        if (_T_563) begin
          if (_T_566) begin
            stateReg <= 4'h9;
          end else begin
            stateReg <= 4'h6;
          end
        end else begin
          stateReg <= 4'ha;
        end
      end else if (_T_503) begin
        stateReg <= 4'h9;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_571) begin
      if (_T_626) begin
        stateReg <= 4'h7;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_628) begin
      if (_T_683) begin
        stateReg <= 4'h8;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_685) begin
      if (_T_502) begin
        stateReg <= 4'h9;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_706) begin
      stateReg <= 4'ha;
    end else if (_T_863) begin
      if (_T_864) begin
        stateReg <= 4'hb;
      end else begin
        stateReg <= 4'hc;
      end
    end else if (_T_887) begin
      stateReg <= 4'hc;
    end else if (_T_978) begin
      stateReg <= 4'hd;
    end else if (_T_1456) begin
      stateReg <= 4'h0;
    end
    if (reset) begin
      shotCnt <= 10'shf;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (!(_T_910)) begin
                                if (!(_T_925)) begin
                                  if (shotPop_0) begin
                                    if (_T_920) begin
                                      shotCnt <= _T_951;
                                    end
                                  end else if (shotPop_1) begin
                                    if (_T_920) begin
                                      shotCnt <= _T_951;
                                    end
                                  end else if (shotPop_2) begin
                                    if (_T_920) begin
                                      shotCnt <= _T_951;
                                    end
                                  end
                                end
                              end
                            end
                          end else if (_T_978) begin
                            if (io_sw_0) begin
                              shotCnt <= 10'shf;
                            end else if (_T_1089) begin
                              if (_T_1100) begin
                                shotCnt <= 10'shf;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      shotLoad <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (_T_910) begin
                                if (shotPop_3) begin
                                  if (_T_920) begin
                                    shotLoad <= 1'h0;
                                  end else begin
                                    shotLoad <= _GEN_887;
                                  end
                                end
                              end else if (_T_925) begin
                                if (shotPop_4) begin
                                  if (_T_920) begin
                                    shotLoad <= 1'h0;
                                  end else begin
                                    shotLoad <= _GEN_902;
                                  end
                                end
                              end else if (shotPop_0) begin
                                if (_T_920) begin
                                  shotLoad <= 1'h0;
                                end else begin
                                  shotLoad <= _GEN_917;
                                end
                              end else if (shotPop_1) begin
                                if (_T_920) begin
                                  shotLoad <= 1'h0;
                                end else begin
                                  shotLoad <= _GEN_917;
                                end
                              end else if (shotPop_2) begin
                                if (_T_920) begin
                                  shotLoad <= 1'h0;
                                end else begin
                                  shotLoad <= _GEN_917;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      shotCntBig <= 3'sh3;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (_T_910) begin
                                if (shotPop_3) begin
                                  if (_T_920) begin
                                    shotCntBig <= _T_923;
                                  end
                                end
                              end
                            end
                          end else if (_T_978) begin
                            if (io_sw_0) begin
                              shotCntBig <= 3'sh3;
                            end else if (_T_1089) begin
                              if (_T_1100) begin
                                shotCntBig <= 3'sh3;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      shotCntFast <= 3'sh3;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (_T_887) begin
                            if (_T_864) begin
                              if (!(_T_910)) begin
                                if (_T_925) begin
                                  if (shotPop_4) begin
                                    if (_T_920) begin
                                      shotCntFast <= _T_938;
                                    end
                                  end
                                end
                              end
                            end
                          end else if (_T_978) begin
                            if (io_sw_0) begin
                              shotCntFast <= 3'sh3;
                            end else if (_T_1089) begin
                              if (_T_1100) begin
                                shotCntFast <= 3'sh3;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    shotPop_0 <= reset | _GEN_4157;
    shotPop_1 <= reset | _GEN_4160;
    shotPop_2 <= reset | _GEN_4163;
    shotPop_3 <= reset | _GEN_4166;
    shotPop_4 <= reset | _GEN_4169;
    shotInteract_0 <= reset | _GEN_4156;
    shotInteract_1 <= reset | _GEN_4159;
    shotInteract_2 <= reset | _GEN_4162;
    shotInteract_3 <= reset | _GEN_4165;
    shotInteract_4 <= reset | _GEN_4168;
    if (reset) begin
      astInteract_0 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_506) begin
      if (_T_508) begin
        if (kill_0_4) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_3) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_2) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_1) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_0) begin
          astInteract_0 <= 1'h0;
        end else if (_T_512) begin
          astInteract_0 <= _GEN_107;
        end else begin
          astInteract_0 <= _GEN_8;
        end
      end else begin
        astInteract_0 <= _GEN_8;
      end
    end else if (_T_571) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_628) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_685) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_0_4) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_3) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_2) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_1) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_0) begin
          astInteract_0 <= 1'h0;
        end else if (_T_512) begin
          astInteract_0 <= _GEN_107;
        end else begin
          astInteract_0 <= _GEN_8;
        end
      end else begin
        astInteract_0 <= _GEN_8;
      end
    end else if (_T_863) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_887) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_978) begin
      if (die_0) begin
        if (_T_1137) begin
          astInteract_0 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_0 <= 1'h0;
        end else begin
          astInteract_0 <= _GEN_8;
        end
      end else if (_T_1086) begin
        astInteract_0 <= 1'h0;
      end else begin
        astInteract_0 <= _GEN_8;
      end
    end else begin
      astInteract_0 <= _GEN_8;
    end
    if (reset) begin
      astInteract_1 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_506) begin
      if (_T_508) begin
        if (kill_1_4) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_3) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_2) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_1) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_0) begin
          astInteract_1 <= 1'h0;
        end else if (_T_512) begin
          astInteract_1 <= _GEN_157;
        end else begin
          astInteract_1 <= _GEN_10;
        end
      end else begin
        astInteract_1 <= _GEN_10;
      end
    end else if (_T_571) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_628) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_685) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_1_4) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_3) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_2) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_1) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_0) begin
          astInteract_1 <= 1'h0;
        end else if (_T_512) begin
          astInteract_1 <= _GEN_157;
        end else begin
          astInteract_1 <= _GEN_10;
        end
      end else begin
        astInteract_1 <= _GEN_10;
      end
    end else if (_T_863) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_887) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_978) begin
      if (die_1) begin
        if (_T_1137) begin
          astInteract_1 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_1 <= 1'h0;
        end else begin
          astInteract_1 <= _GEN_10;
        end
      end else if (_T_1086) begin
        astInteract_1 <= 1'h0;
      end else begin
        astInteract_1 <= _GEN_10;
      end
    end else begin
      astInteract_1 <= _GEN_10;
    end
    if (reset) begin
      astInteract_2 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_506) begin
      if (_T_508) begin
        if (kill_2_4) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_3) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_2) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_1) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_0) begin
          astInteract_2 <= 1'h0;
        end else if (_T_512) begin
          astInteract_2 <= _GEN_207;
        end else begin
          astInteract_2 <= _GEN_12;
        end
      end else begin
        astInteract_2 <= _GEN_12;
      end
    end else if (_T_571) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_628) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_685) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_2_4) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_3) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_2) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_1) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_0) begin
          astInteract_2 <= 1'h0;
        end else if (_T_512) begin
          astInteract_2 <= _GEN_207;
        end else begin
          astInteract_2 <= _GEN_12;
        end
      end else begin
        astInteract_2 <= _GEN_12;
      end
    end else if (_T_863) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_887) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_978) begin
      if (die_2) begin
        if (_T_1137) begin
          astInteract_2 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_2 <= 1'h0;
        end else begin
          astInteract_2 <= _GEN_12;
        end
      end else if (_T_1086) begin
        astInteract_2 <= 1'h0;
      end else begin
        astInteract_2 <= _GEN_12;
      end
    end else begin
      astInteract_2 <= _GEN_12;
    end
    if (reset) begin
      astInteract_3 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_506) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_571) begin
      if (kill_3_4) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_3) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_2) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_1) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_0) begin
        astInteract_3 <= 1'h0;
      end else if (_T_512) begin
        astInteract_3 <= _GEN_285;
      end else begin
        astInteract_3 <= _GEN_14;
      end
    end else if (_T_628) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_685) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_706) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_863) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_887) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_978) begin
      if (die_3) begin
        if (_T_1137) begin
          astInteract_3 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_3 <= 1'h0;
        end else begin
          astInteract_3 <= _GEN_14;
        end
      end else if (_T_1086) begin
        astInteract_3 <= 1'h0;
      end else begin
        astInteract_3 <= _GEN_14;
      end
    end else begin
      astInteract_3 <= _GEN_14;
    end
    if (reset) begin
      astInteract_4 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_506) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_571) begin
      if (kill_4_4) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_3) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_2) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_1) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_0) begin
        astInteract_4 <= 1'h0;
      end else if (_T_512) begin
        astInteract_4 <= _GEN_335;
      end else begin
        astInteract_4 <= _GEN_16;
      end
    end else if (_T_628) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_685) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_4_4) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_3) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_2) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_1) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_0) begin
          astInteract_4 <= 1'h0;
        end else if (_T_512) begin
          astInteract_4 <= _GEN_335;
        end else begin
          astInteract_4 <= _GEN_16;
        end
      end else begin
        astInteract_4 <= _GEN_16;
      end
    end else if (_T_863) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_887) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_978) begin
      if (die_4) begin
        if (_T_1137) begin
          astInteract_4 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_4 <= 1'h0;
        end else begin
          astInteract_4 <= _GEN_16;
        end
      end else if (_T_1086) begin
        astInteract_4 <= 1'h0;
      end else begin
        astInteract_4 <= _GEN_16;
      end
    end else begin
      astInteract_4 <= _GEN_16;
    end
    if (reset) begin
      astInteract_5 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_506) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_571) begin
      if (kill_5_4) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_3) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_2) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_1) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_0) begin
        astInteract_5 <= 1'h0;
      end else if (_T_512) begin
        astInteract_5 <= _GEN_385;
      end else begin
        astInteract_5 <= _GEN_18;
      end
    end else if (_T_628) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_685) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_5_4) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_3) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_2) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_1) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_0) begin
          astInteract_5 <= 1'h0;
        end else if (_T_512) begin
          astInteract_5 <= _GEN_385;
        end else begin
          astInteract_5 <= _GEN_18;
        end
      end else begin
        astInteract_5 <= _GEN_18;
      end
    end else if (_T_863) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_887) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_978) begin
      if (die_5) begin
        if (_T_1137) begin
          astInteract_5 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_5 <= 1'h0;
        end else begin
          astInteract_5 <= _GEN_18;
        end
      end else if (_T_1086) begin
        astInteract_5 <= 1'h0;
      end else begin
        astInteract_5 <= _GEN_18;
      end
    end else begin
      astInteract_5 <= _GEN_18;
    end
    if (reset) begin
      astInteract_6 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_506) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_571) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_628) begin
      if (kill_6_4) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_3) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_2) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_1) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_0) begin
        astInteract_6 <= 1'h0;
      end else if (_T_512) begin
        astInteract_6 <= _GEN_435;
      end else begin
        astInteract_6 <= _GEN_20;
      end
    end else if (_T_685) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_706) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_863) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_887) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_978) begin
      if (die_6) begin
        if (_T_1137) begin
          astInteract_6 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_6 <= 1'h0;
        end else begin
          astInteract_6 <= _GEN_20;
        end
      end else if (_T_1086) begin
        astInteract_6 <= 1'h0;
      end else begin
        astInteract_6 <= _GEN_20;
      end
    end else begin
      astInteract_6 <= _GEN_20;
    end
    if (reset) begin
      astInteract_7 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_506) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_571) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_628) begin
      if (kill_7_4) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_3) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_2) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_1) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_0) begin
        astInteract_7 <= 1'h0;
      end else if (_T_512) begin
        astInteract_7 <= _GEN_485;
      end else begin
        astInteract_7 <= _GEN_22;
      end
    end else if (_T_685) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_706) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_863) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_887) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_978) begin
      if (die_7) begin
        if (_T_1137) begin
          astInteract_7 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_7 <= 1'h0;
        end else begin
          astInteract_7 <= _GEN_22;
        end
      end else if (_T_1086) begin
        astInteract_7 <= 1'h0;
      end else begin
        astInteract_7 <= _GEN_22;
      end
    end else begin
      astInteract_7 <= _GEN_22;
    end
    if (reset) begin
      astInteract_8 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_506) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_571) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_628) begin
      if (kill_8_4) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_3) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_2) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_1) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_0) begin
        astInteract_8 <= 1'h0;
      end else if (_T_512) begin
        astInteract_8 <= _GEN_535;
      end else begin
        astInteract_8 <= _GEN_24;
      end
    end else if (_T_685) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_706) begin
      astInteract_8 <= 1'h0;
    end else if (_T_863) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_887) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_978) begin
      if (die_8) begin
        if (_T_1137) begin
          astInteract_8 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_8 <= 1'h0;
        end else begin
          astInteract_8 <= _GEN_24;
        end
      end else if (_T_1086) begin
        astInteract_8 <= 1'h0;
      end else begin
        astInteract_8 <= _GEN_24;
      end
    end else begin
      astInteract_8 <= _GEN_24;
    end
    if (reset) begin
      astInteract_9 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_506) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_571) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_628) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_685) begin
      if (kill_9_3) begin
        astInteract_9 <= 1'h0;
      end else if (_T_689) begin
        astInteract_9 <= _GEN_585;
      end else begin
        astInteract_9 <= _GEN_26;
      end
    end else if (_T_706) begin
      if (_T_707) begin
        if (kill_9_3) begin
          astInteract_9 <= 1'h0;
        end else if (_T_689) begin
          astInteract_9 <= _GEN_585;
        end else begin
          astInteract_9 <= _GEN_26;
        end
      end else begin
        astInteract_9 <= _GEN_26;
      end
    end else if (_T_863) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_887) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_978) begin
      if (die_9) begin
        if (_T_1137) begin
          astInteract_9 <= 1'h0;
        end else if (_T_1086) begin
          astInteract_9 <= 1'h0;
        end else begin
          astInteract_9 <= _GEN_26;
        end
      end else if (_T_1086) begin
        astInteract_9 <= 1'h0;
      end else begin
        astInteract_9 <= _GEN_26;
      end
    end else begin
      astInteract_9 <= _GEN_26;
    end
    if (reset) begin
      astInteract_10 <= 1'h0;
    end else if (_T_342) begin
      if (_T_341) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_343) begin
      if (_T_341) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_405) begin
      if (_T_341) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_452) begin
      if (_T_341) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_487) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_506) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_571) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_628) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_685) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_706) begin
      if (_T_501) begin
        astInteract_10 <= 1'h0;
      end else if (_T_831) begin
        astInteract_10 <= _GEN_826;
      end else begin
        astInteract_10 <= _GEN_28;
      end
    end else if (_T_863) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_887) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_978) begin
      if (die_10) begin
        if (_T_1137) begin
          astInteract_10 <= 1'h0;
        end else begin
          astInteract_10 <= _GEN_28;
        end
      end else begin
        astInteract_10 <= _GEN_28;
      end
    end else begin
      astInteract_10 <= _GEN_28;
    end
    shipInteract <= reset | _GEN_4255;
    if (reset) begin
      die_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_0 <= _T_1124;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_1 <= _T_1141;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_2 <= _T_1158;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_3 <= _T_1175;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_4 <= _T_1192;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_5 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_5 <= _T_1209;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_6 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_6 <= _T_1226;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_7 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_7 <= _T_1243;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_8 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_8 <= _T_1260;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_9 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_9 <= _T_1277;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_10 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              die_10 <= _T_1294;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_0_0 <= _T_1126;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_0_1 <= _T_1128;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_0_2 <= _T_1130;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_0_3 <= _T_1132;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_0_4 <= _T_1134;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_1_0 <= _T_1143;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_1_1 <= _T_1145;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_1_2 <= _T_1147;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_1_3 <= _T_1149;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_1_4 <= _T_1151;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_2_0 <= _T_1160;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_2_1 <= _T_1162;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_2_2 <= _T_1164;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_2_3 <= _T_1166;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_2_4 <= _T_1168;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_3_0 <= _T_1177;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_3_1 <= _T_1179;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_3_2 <= _T_1181;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_3_3 <= _T_1183;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_3_4 <= _T_1185;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_4_0 <= _T_1194;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_4_1 <= _T_1196;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_4_2 <= _T_1198;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_4_3 <= _T_1200;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_4_4 <= _T_1202;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_5_0 <= _T_1211;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_5_1 <= _T_1213;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_5_2 <= _T_1215;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_5_3 <= _T_1217;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_5_4 <= _T_1219;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_6_0 <= _T_1228;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_6_1 <= _T_1230;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_6_2 <= _T_1232;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_6_3 <= _T_1234;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_6_4 <= _T_1236;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_7_0 <= _T_1245;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_7_1 <= _T_1247;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_7_2 <= _T_1249;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_7_3 <= _T_1251;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_7_4 <= _T_1253;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_8_0 <= _T_1262;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_8_1 <= _T_1264;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_8_2 <= _T_1266;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_8_3 <= _T_1268;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_8_4 <= _T_1270;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_9_0 <= _T_1279;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_9_1 <= _T_1281;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_9_2 <= _T_1283;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_9_3 <= _T_1285;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_0 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_10_0 <= _T_1296;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_1 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_10_1 <= _T_1298;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_2 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_10_2 <= _T_1300;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_3 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_10_3 <= _T_1302;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_4 <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              kill_10_4 <= _T_1304;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      hp <= 4'h3;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (io_sw_0) begin
                                hp <= 4'h3;
                              end else if (die_10) begin
                                if (_T_1137) begin
                                  hp <= _T_1139;
                                end else if (die_9) begin
                                  if (_T_1137) begin
                                    hp <= _T_1139;
                                  end else if (die_8) begin
                                    if (_T_1137) begin
                                      hp <= _T_1139;
                                    end else if (die_7) begin
                                      if (_T_1137) begin
                                        hp <= _T_1139;
                                      end else if (die_6) begin
                                        if (_T_1137) begin
                                          hp <= _T_1139;
                                        end else if (die_5) begin
                                          if (_T_1137) begin
                                            hp <= _T_1139;
                                          end else if (die_4) begin
                                            if (_T_1137) begin
                                              hp <= _T_1139;
                                            end else if (die_3) begin
                                              if (_T_1137) begin
                                                hp <= _T_1139;
                                              end else if (die_2) begin
                                                if (_T_1137) begin
                                                  hp <= _T_1139;
                                                end else if (die_1) begin
                                                  if (_T_1137) begin
                                                    hp <= _T_1139;
                                                  end else if (die_0) begin
                                                    if (_T_1137) begin
                                                      hp <= _T_1139;
                                                    end else if (_T_1089) begin
                                                      if (_T_1100) begin
                                                        hp <= 4'h3;
                                                      end
                                                    end
                                                  end else if (_T_1089) begin
                                                    if (_T_1100) begin
                                                      hp <= 4'h3;
                                                    end
                                                  end
                                                end else if (die_0) begin
                                                  if (_T_1137) begin
                                                    hp <= _T_1139;
                                                  end else if (_T_1089) begin
                                                    if (_T_1100) begin
                                                      hp <= 4'h3;
                                                    end
                                                  end
                                                end else if (_T_1089) begin
                                                  if (_T_1100) begin
                                                    hp <= 4'h3;
                                                  end
                                                end
                                              end else if (die_1) begin
                                                if (_T_1137) begin
                                                  hp <= _T_1139;
                                                end else if (die_0) begin
                                                  if (_T_1137) begin
                                                    hp <= _T_1139;
                                                  end else begin
                                                    hp <= _GEN_1169;
                                                  end
                                                end else begin
                                                  hp <= _GEN_1169;
                                                end
                                              end else if (die_0) begin
                                                if (_T_1137) begin
                                                  hp <= _T_1139;
                                                end else begin
                                                  hp <= _GEN_1169;
                                                end
                                              end else begin
                                                hp <= _GEN_1169;
                                              end
                                            end else if (die_2) begin
                                              if (_T_1137) begin
                                                hp <= _T_1139;
                                              end else if (die_1) begin
                                                if (_T_1137) begin
                                                  hp <= _T_1139;
                                                end else begin
                                                  hp <= _GEN_1184;
                                                end
                                              end else begin
                                                hp <= _GEN_1184;
                                              end
                                            end else if (die_1) begin
                                              if (_T_1137) begin
                                                hp <= _T_1139;
                                              end else begin
                                                hp <= _GEN_1184;
                                              end
                                            end else begin
                                              hp <= _GEN_1184;
                                            end
                                          end else if (die_3) begin
                                            if (_T_1137) begin
                                              hp <= _T_1139;
                                            end else if (die_2) begin
                                              if (_T_1137) begin
                                                hp <= _T_1139;
                                              end else begin
                                                hp <= _GEN_1194;
                                              end
                                            end else begin
                                              hp <= _GEN_1194;
                                            end
                                          end else if (die_2) begin
                                            if (_T_1137) begin
                                              hp <= _T_1139;
                                            end else begin
                                              hp <= _GEN_1194;
                                            end
                                          end else begin
                                            hp <= _GEN_1194;
                                          end
                                        end else if (die_4) begin
                                          if (_T_1137) begin
                                            hp <= _T_1139;
                                          end else if (die_3) begin
                                            if (_T_1137) begin
                                              hp <= _T_1139;
                                            end else begin
                                              hp <= _GEN_1204;
                                            end
                                          end else begin
                                            hp <= _GEN_1204;
                                          end
                                        end else if (die_3) begin
                                          if (_T_1137) begin
                                            hp <= _T_1139;
                                          end else begin
                                            hp <= _GEN_1204;
                                          end
                                        end else begin
                                          hp <= _GEN_1204;
                                        end
                                      end else if (die_5) begin
                                        if (_T_1137) begin
                                          hp <= _T_1139;
                                        end else if (die_4) begin
                                          if (_T_1137) begin
                                            hp <= _T_1139;
                                          end else begin
                                            hp <= _GEN_1214;
                                          end
                                        end else begin
                                          hp <= _GEN_1214;
                                        end
                                      end else if (die_4) begin
                                        if (_T_1137) begin
                                          hp <= _T_1139;
                                        end else begin
                                          hp <= _GEN_1214;
                                        end
                                      end else begin
                                        hp <= _GEN_1214;
                                      end
                                    end else if (die_6) begin
                                      if (_T_1137) begin
                                        hp <= _T_1139;
                                      end else if (die_5) begin
                                        if (_T_1137) begin
                                          hp <= _T_1139;
                                        end else begin
                                          hp <= _GEN_1224;
                                        end
                                      end else begin
                                        hp <= _GEN_1224;
                                      end
                                    end else if (die_5) begin
                                      if (_T_1137) begin
                                        hp <= _T_1139;
                                      end else begin
                                        hp <= _GEN_1224;
                                      end
                                    end else begin
                                      hp <= _GEN_1224;
                                    end
                                  end else if (die_7) begin
                                    if (_T_1137) begin
                                      hp <= _T_1139;
                                    end else if (die_6) begin
                                      if (_T_1137) begin
                                        hp <= _T_1139;
                                      end else begin
                                        hp <= _GEN_1234;
                                      end
                                    end else begin
                                      hp <= _GEN_1234;
                                    end
                                  end else if (die_6) begin
                                    if (_T_1137) begin
                                      hp <= _T_1139;
                                    end else begin
                                      hp <= _GEN_1234;
                                    end
                                  end else begin
                                    hp <= _GEN_1234;
                                  end
                                end else if (die_8) begin
                                  if (_T_1137) begin
                                    hp <= _T_1139;
                                  end else if (die_7) begin
                                    if (_T_1137) begin
                                      hp <= _T_1139;
                                    end else begin
                                      hp <= _GEN_1244;
                                    end
                                  end else begin
                                    hp <= _GEN_1244;
                                  end
                                end else if (die_7) begin
                                  if (_T_1137) begin
                                    hp <= _T_1139;
                                  end else begin
                                    hp <= _GEN_1244;
                                  end
                                end else begin
                                  hp <= _GEN_1244;
                                end
                              end else if (die_9) begin
                                if (_T_1137) begin
                                  hp <= _T_1139;
                                end else if (die_8) begin
                                  if (_T_1137) begin
                                    hp <= _T_1139;
                                  end else begin
                                    hp <= _GEN_1254;
                                  end
                                end else begin
                                  hp <= _GEN_1254;
                                end
                              end else if (die_8) begin
                                if (_T_1137) begin
                                  hp <= _T_1139;
                                end else begin
                                  hp <= _GEN_1254;
                                end
                              end else begin
                                hp <= _GEN_1254;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      planetHp <= 5'ha;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (_T_706) begin
                        if (kill_10_4) begin
                          if (_T_689) begin
                            planetHp <= _T_849;
                          end else if (kill_10_3) begin
                            if (_T_689) begin
                              planetHp <= _T_849;
                            end else if (kill_10_2) begin
                              if (_T_689) begin
                                planetHp <= _T_849;
                              end else if (kill_10_1) begin
                                if (_T_689) begin
                                  planetHp <= _T_849;
                                end else if (kill_10_0) begin
                                  if (_T_689) begin
                                    planetHp <= _T_849;
                                  end
                                end
                              end else if (kill_10_0) begin
                                if (_T_689) begin
                                  planetHp <= _T_849;
                                end
                              end
                            end else if (kill_10_1) begin
                              if (_T_689) begin
                                planetHp <= _T_849;
                              end else if (kill_10_0) begin
                                if (_T_689) begin
                                  planetHp <= _T_849;
                                end
                              end
                            end else if (kill_10_0) begin
                              if (_T_689) begin
                                planetHp <= _T_849;
                              end
                            end
                          end else if (kill_10_2) begin
                            if (_T_689) begin
                              planetHp <= _T_849;
                            end else if (kill_10_1) begin
                              if (_T_689) begin
                                planetHp <= _T_849;
                              end else begin
                                planetHp <= _GEN_835;
                              end
                            end else begin
                              planetHp <= _GEN_835;
                            end
                          end else if (kill_10_1) begin
                            if (_T_689) begin
                              planetHp <= _T_849;
                            end else begin
                              planetHp <= _GEN_835;
                            end
                          end else begin
                            planetHp <= _GEN_835;
                          end
                        end else if (kill_10_3) begin
                          if (_T_689) begin
                            planetHp <= _T_849;
                          end else if (kill_10_2) begin
                            if (_T_689) begin
                              planetHp <= _T_849;
                            end else begin
                              planetHp <= _GEN_840;
                            end
                          end else begin
                            planetHp <= _GEN_840;
                          end
                        end else if (kill_10_2) begin
                          if (_T_689) begin
                            planetHp <= _T_849;
                          end else begin
                            planetHp <= _GEN_840;
                          end
                        end else begin
                          planetHp <= _GEN_840;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spwnProt <= 6'sh0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1315) begin
                                spwnProt <= 6'sh0;
                              end else if (_T_1311) begin
                                spwnProt <= _T_1314;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    show <= reset | _GEN_4246;
    if (reset) begin
      blink <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              blink <= _T_1117;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      secCnt <= 8'sh0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1089) begin
                                if (_T_1100) begin
                                  secCnt <= 8'sh0;
                                end else if (_T_1105) begin
                                  secCnt <= 8'shf;
                                end else begin
                                  secCnt <= _T_1092;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      level <= 3'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1089) begin
                                if (_T_1100) begin
                                  level <= _T_1102;
                                end else if (_T_501) begin
                                  level <= 3'h5;
                                end
                              end else if (_T_501) begin
                                level <= 3'h5;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      start <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              start <= _GEN_1294;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      levelCng <= 1'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (_T_405) begin
          if (_T_406) begin
            levelCng <= 1'h0;
          end
        end else if (!(_T_452)) begin
          if (!(_T_487)) begin
            if (!(_T_506)) begin
              if (!(_T_571)) begin
                if (!(_T_628)) begin
                  if (!(_T_685)) begin
                    if (!(_T_706)) begin
                      if (!(_T_863)) begin
                        if (!(_T_887)) begin
                          if (_T_978) begin
                            if (_T_1089) begin
                              levelCng <= _GEN_1167;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cngCnt <= 4'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1119) begin
                                if (_T_1122) begin
                                  cngCnt <= 4'h0;
                                end else begin
                                  cngCnt <= _T_1121;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cnt <= 10'sh0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1088) begin
                                cnt <= 10'sh0;
                              end else begin
                                cnt <= _T_1109;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      count1 <= 7'h0;
    end else if (!(_T_342)) begin
      if (_T_343) begin
        if (_T_396) begin
          if (levelCng) begin
            count1 <= _T_404;
          end
        end
      end else if (_T_405) begin
        if (_T_406) begin
          count1 <= 7'h0;
        end
      end else if (_T_452) begin
        if (_T_407) begin
          if (_T_408) begin
            count1 <= _T_404;
          end
        end
      end
    end
    if (reset) begin
      count3 <= 7'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (_T_405) begin
          if (_T_438) begin
            if (_T_409) begin
              count3 <= _T_421;
            end else begin
              count3 <= 7'h0;
            end
          end else if (_T_424) begin
            if (_T_409) begin
              count3 <= _T_421;
            end else begin
              count3 <= 7'h0;
            end
          end else if (_T_407) begin
            if (_T_408) begin
              if (_T_409) begin
                count3 <= _T_421;
              end else begin
                count3 <= 7'h0;
              end
            end
          end
        end else if (_T_452) begin
          if (_T_438) begin
            if (_T_409) begin
              count3 <= _T_421;
            end else begin
              count3 <= 7'h0;
            end
          end else if (_T_424) begin
            count3 <= _GEN_40;
          end
        end else if (_T_487) begin
          if (_T_409) begin
            count3 <= _T_421;
          end else if (!(_T_501)) begin
            count3 <= 7'h0;
          end
        end
      end
    end
    if (reset) begin
      count4 <= 8'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (_T_452) begin
            if (_T_424) begin
              if (_T_409) begin
                if (_T_407) begin
                  if (_T_408) begin
                    count4 <= 8'h0;
                  end
                end
              end else begin
                count4 <= 8'h1;
              end
            end else if (_T_407) begin
              if (_T_408) begin
                count4 <= 8'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      count5 <= 8'h0;
    end else if (!(_T_342)) begin
      if (!(_T_343)) begin
        if (!(_T_405)) begin
          if (!(_T_452)) begin
            if (!(_T_487)) begin
              if (!(_T_506)) begin
                if (!(_T_571)) begin
                  if (!(_T_628)) begin
                    if (!(_T_685)) begin
                      if (!(_T_706)) begin
                        if (!(_T_863)) begin
                          if (!(_T_887)) begin
                            if (_T_978) begin
                              if (_T_1027) begin
                                count5 <= 8'h1;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    _T_913 <= Xstart_0;
    _T_918 <= Ystart_0;
    _T_928 <= Xstart_0;
    _T_933 <= Ystart_0;
    _T_941 <= Xstart_0;
    _T_946 <= Ystart_0;
    _T_954 <= Xstart_0;
    _T_959 <= Ystart_0;
    _T_967 <= Xstart_0;
    _T_972 <= Ystart_0;
    if (reset) begin
      _T_979 <= 1'h0;
    end else begin
      _T_979 <= _GEN_1078;
    end
    if (reset) begin
      _T_980 <= 1'h0;
    end else begin
      _T_980 <= _GEN_1079;
    end
    if (reset) begin
      _T_981 <= 3'sh0;
    end else if (_T_984) begin
      _T_981 <= {{1{Randomizer_33_io_out[1]}},Randomizer_33_io_out};
    end
    if (reset) begin
      _T_982 <= 3'sh0;
    end else if (_T_985) begin
      _T_982 <= {{1{Randomizer_33_io_out[1]}},Randomizer_33_io_out};
    end
    if (reset) begin
      _T_983 <= 3'sh0;
    end else if (_T_986) begin
      _T_983 <= {{1{Randomizer_33_io_out[1]}},Randomizer_33_io_out};
    end
    if (reset) begin
      _T_1029 <= 1'h0;
    end else begin
      _T_1029 <= _GEN_1107;
    end
    if (reset) begin
      _T_1030 <= 1'h0;
    end else begin
      _T_1030 <= _GEN_1108;
    end
    if (reset) begin
      _T_1031 <= 3'sh0;
    end else if (_T_1034) begin
      _T_1031 <= {{1{Randomizer_40_io_out[1]}},Randomizer_40_io_out};
    end
    if (reset) begin
      _T_1032 <= 3'sh0;
    end else if (_T_1035) begin
      _T_1032 <= {{1{Randomizer_40_io_out[1]}},Randomizer_40_io_out};
    end
    if (reset) begin
      _T_1033 <= 3'sh0;
    end else if (_T_1036) begin
      _T_1033 <= {{1{Randomizer_40_io_out[1]}},Randomizer_40_io_out};
    end
  end
endmodule
module GameTop(
  input        clock,
  input        reset,
  input        io_btnC,
  input        io_btnU,
  input        io_btnL,
  input        io_btnR,
  input        io_btnD,
  output [3:0] io_vgaRed,
  output [3:0] io_vgaBlue,
  output [3:0] io_vgaGreen,
  output       io_Hsync,
  output       io_Vsync,
  input        io_sw_0,
  input        io_sw_1,
  input        io_sw_2,
  input        io_sw_7,
  output       io_soundOutput_0,
  output       io_missingFrameError,
  output       io_backBufferWriteError,
  output       io_viewBoxOutOfRangeError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire  graphicEngineVGA_clock; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_reset; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_0; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_1; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_2; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_3; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_4; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_5; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_6; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_7; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_8; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_9; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_10; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_11; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_12; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_13; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_14; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_15; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_16; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_17; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_18; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_19; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_20; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_21; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_22; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_23; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_24; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_25; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_26; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_27; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_28; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_29; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_30; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_31; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_32; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_33; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_41; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_42; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_43; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_44; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_45; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_46; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_47; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_48; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_49; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_50; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_51; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_122; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_123; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_124; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_125; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_126; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_127; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_0; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_1; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_2; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_3; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_4; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_5; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_6; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_7; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_8; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_9; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_10; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_11; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_12; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_13; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_14; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_15; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_16; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_17; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_18; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_19; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_20; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_21; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_22; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_23; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_24; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_25; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_26; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_27; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_28; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_29; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_30; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_31; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_32; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_33; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_41; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_42; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_43; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_122; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_123; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_124; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_125; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_126; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_127; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_0; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_1; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_2; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_3; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_4; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_5; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_6; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_7; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_8; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_9; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_10; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_11; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_12; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_13; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_14; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_15; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_16; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_17; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_18; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_19; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_20; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_21; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_22; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_23; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_24; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_25; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_26; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_27; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_28; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_29; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_30; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_31; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_32; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_33; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_41; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_42; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_43; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_44; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_45; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_46; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_47; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_48; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_49; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_50; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_51; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_55; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_56; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_57; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_61; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_62; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_63; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_64; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_65; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_66; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_70; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_71; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_72; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_122; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_123; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_124; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_125; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_126; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_127; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_viewBoxX_0; // @[GameTop.scala 46:32]
  wire [4:0] graphicEngineVGA_io_backBufferWriteData; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_backBufferWriteAddress; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_backBufferWriteEnable; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_newFrame; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_frameUpdateDone; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_missingFrameError; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_backBufferWriteError; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_viewBoxOutOfRangeError; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaRed; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaBlue; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaGreen; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Hsync; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Vsync; // @[GameTop.scala 46:32]
  wire  soundEngine_clock; // @[GameTop.scala 48:27]
  wire  soundEngine_reset; // @[GameTop.scala 48:27]
  wire  soundEngine_io_output_0; // @[GameTop.scala 48:27]
  wire [3:0] soundEngine_io_input; // @[GameTop.scala 48:27]
  wire  gameLogic_clock; // @[GameTop.scala 52:25]
  wire  gameLogic_reset; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnC; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnU; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnL; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnR; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnD; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_0; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_1; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_2; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_7; // @[GameTop.scala 52:25]
  wire [3:0] gameLogic_io_songInput; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_0; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_1; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_2; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_3; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_4; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_5; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_6; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_7; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_8; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_9; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_10; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_11; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_12; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_13; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_14; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_15; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_16; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_17; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_18; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_19; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_20; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_21; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_22; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_23; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_24; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_25; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_26; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_27; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_28; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_29; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_30; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_31; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_32; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_33; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_41; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_42; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_43; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_44; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_45; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_46; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_47; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_48; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_49; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_50; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_51; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_122; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_123; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_124; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_125; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_126; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_127; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_0; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_1; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_2; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_3; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_4; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_5; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_6; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_7; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_8; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_9; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_10; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_11; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_12; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_13; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_14; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_15; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_16; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_17; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_18; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_19; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_20; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_21; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_22; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_23; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_24; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_25; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_26; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_27; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_28; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_29; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_30; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_31; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_32; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_33; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_41; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_42; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_43; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_122; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_123; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_124; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_125; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_126; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_127; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_0; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_1; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_2; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_3; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_4; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_5; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_6; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_7; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_8; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_9; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_10; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_11; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_12; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_13; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_14; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_15; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_16; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_17; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_18; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_19; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_20; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_21; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_22; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_23; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_24; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_25; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_26; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_27; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_28; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_29; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_30; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_31; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_32; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_33; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_41; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_42; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_43; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_44; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_45; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_46; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_47; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_48; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_49; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_50; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_51; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_55; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_56; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_57; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_61; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_62; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_63; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_64; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_65; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_66; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_70; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_71; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_72; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_122; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_123; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_124; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_125; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_126; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_127; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_viewBoxX_0; // @[GameTop.scala 52:25]
  wire [4:0] gameLogic_io_backBufferWriteData; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_backBufferWriteAddress; // @[GameTop.scala 52:25]
  wire  gameLogic_io_backBufferWriteEnable; // @[GameTop.scala 52:25]
  wire  gameLogic_io_newFrame; // @[GameTop.scala 52:25]
  wire  gameLogic_io_frameUpdateDone; // @[GameTop.scala 52:25]
  reg [20:0] debounceCounter; // @[GameTop.scala 73:32]
  wire  debounceSampleEn = debounceCounter == 21'h1e847f; // @[GameTop.scala 75:24]
  wire [20:0] _T_2 = debounceCounter + 21'h1; // @[GameTop.scala 79:40]
  reg [21:0] resetReleaseCounter; // @[GameTop.scala 86:36]
  wire  _T_3 = resetReleaseCounter == 22'h3d08ff; // @[GameTop.scala 88:28]
  wire [21:0] _T_5 = resetReleaseCounter + 22'h1; // @[GameTop.scala 92:48]
  reg  _T_7_0; // @[GameUtilities.scala 39:28]
  reg  _T_7_1; // @[GameUtilities.scala 39:28]
  reg  _T_7_2; // @[GameUtilities.scala 39:28]
  reg  btnCState; // @[Reg.scala 27:20]
  reg  _T_9_0; // @[GameUtilities.scala 39:28]
  reg  _T_9_1; // @[GameUtilities.scala 39:28]
  reg  _T_9_2; // @[GameUtilities.scala 39:28]
  reg  btnUState; // @[Reg.scala 27:20]
  reg  _T_11_0; // @[GameUtilities.scala 39:28]
  reg  _T_11_1; // @[GameUtilities.scala 39:28]
  reg  _T_11_2; // @[GameUtilities.scala 39:28]
  reg  btnLState; // @[Reg.scala 27:20]
  reg  _T_13_0; // @[GameUtilities.scala 39:28]
  reg  _T_13_1; // @[GameUtilities.scala 39:28]
  reg  _T_13_2; // @[GameUtilities.scala 39:28]
  reg  btnRState; // @[Reg.scala 27:20]
  reg  _T_15_0; // @[GameUtilities.scala 39:28]
  reg  _T_15_1; // @[GameUtilities.scala 39:28]
  reg  _T_15_2; // @[GameUtilities.scala 39:28]
  reg  btnDState; // @[Reg.scala 27:20]
  reg  _T_17_0; // @[GameUtilities.scala 39:28]
  reg  _T_17_1; // @[GameUtilities.scala 39:28]
  reg  _T_17_2; // @[GameUtilities.scala 39:28]
  reg  _T_18; // @[Reg.scala 27:20]
  reg  _T_20_0; // @[GameUtilities.scala 39:28]
  reg  _T_20_1; // @[GameUtilities.scala 39:28]
  reg  _T_20_2; // @[GameUtilities.scala 39:28]
  reg  _T_21; // @[Reg.scala 27:20]
  reg  _T_23_0; // @[GameUtilities.scala 39:28]
  reg  _T_23_1; // @[GameUtilities.scala 39:28]
  reg  _T_23_2; // @[GameUtilities.scala 39:28]
  reg  _T_24; // @[Reg.scala 27:20]
  reg  _T_38_0; // @[GameUtilities.scala 39:28]
  reg  _T_38_1; // @[GameUtilities.scala 39:28]
  reg  _T_38_2; // @[GameUtilities.scala 39:28]
  reg  _T_39; // @[Reg.scala 27:20]
  GraphicEngineVGA graphicEngineVGA ( // @[GameTop.scala 46:32]
    .clock(graphicEngineVGA_clock),
    .reset(graphicEngineVGA_reset),
    .io_spriteXPosition_0(graphicEngineVGA_io_spriteXPosition_0),
    .io_spriteXPosition_1(graphicEngineVGA_io_spriteXPosition_1),
    .io_spriteXPosition_2(graphicEngineVGA_io_spriteXPosition_2),
    .io_spriteXPosition_3(graphicEngineVGA_io_spriteXPosition_3),
    .io_spriteXPosition_4(graphicEngineVGA_io_spriteXPosition_4),
    .io_spriteXPosition_5(graphicEngineVGA_io_spriteXPosition_5),
    .io_spriteXPosition_6(graphicEngineVGA_io_spriteXPosition_6),
    .io_spriteXPosition_7(graphicEngineVGA_io_spriteXPosition_7),
    .io_spriteXPosition_8(graphicEngineVGA_io_spriteXPosition_8),
    .io_spriteXPosition_9(graphicEngineVGA_io_spriteXPosition_9),
    .io_spriteXPosition_10(graphicEngineVGA_io_spriteXPosition_10),
    .io_spriteXPosition_11(graphicEngineVGA_io_spriteXPosition_11),
    .io_spriteXPosition_12(graphicEngineVGA_io_spriteXPosition_12),
    .io_spriteXPosition_13(graphicEngineVGA_io_spriteXPosition_13),
    .io_spriteXPosition_14(graphicEngineVGA_io_spriteXPosition_14),
    .io_spriteXPosition_15(graphicEngineVGA_io_spriteXPosition_15),
    .io_spriteXPosition_16(graphicEngineVGA_io_spriteXPosition_16),
    .io_spriteXPosition_17(graphicEngineVGA_io_spriteXPosition_17),
    .io_spriteXPosition_18(graphicEngineVGA_io_spriteXPosition_18),
    .io_spriteXPosition_19(graphicEngineVGA_io_spriteXPosition_19),
    .io_spriteXPosition_20(graphicEngineVGA_io_spriteXPosition_20),
    .io_spriteXPosition_21(graphicEngineVGA_io_spriteXPosition_21),
    .io_spriteXPosition_22(graphicEngineVGA_io_spriteXPosition_22),
    .io_spriteXPosition_23(graphicEngineVGA_io_spriteXPosition_23),
    .io_spriteXPosition_24(graphicEngineVGA_io_spriteXPosition_24),
    .io_spriteXPosition_25(graphicEngineVGA_io_spriteXPosition_25),
    .io_spriteXPosition_26(graphicEngineVGA_io_spriteXPosition_26),
    .io_spriteXPosition_27(graphicEngineVGA_io_spriteXPosition_27),
    .io_spriteXPosition_28(graphicEngineVGA_io_spriteXPosition_28),
    .io_spriteXPosition_29(graphicEngineVGA_io_spriteXPosition_29),
    .io_spriteXPosition_30(graphicEngineVGA_io_spriteXPosition_30),
    .io_spriteXPosition_31(graphicEngineVGA_io_spriteXPosition_31),
    .io_spriteXPosition_32(graphicEngineVGA_io_spriteXPosition_32),
    .io_spriteXPosition_33(graphicEngineVGA_io_spriteXPosition_33),
    .io_spriteXPosition_41(graphicEngineVGA_io_spriteXPosition_41),
    .io_spriteXPosition_42(graphicEngineVGA_io_spriteXPosition_42),
    .io_spriteXPosition_43(graphicEngineVGA_io_spriteXPosition_43),
    .io_spriteXPosition_44(graphicEngineVGA_io_spriteXPosition_44),
    .io_spriteXPosition_45(graphicEngineVGA_io_spriteXPosition_45),
    .io_spriteXPosition_46(graphicEngineVGA_io_spriteXPosition_46),
    .io_spriteXPosition_47(graphicEngineVGA_io_spriteXPosition_47),
    .io_spriteXPosition_48(graphicEngineVGA_io_spriteXPosition_48),
    .io_spriteXPosition_49(graphicEngineVGA_io_spriteXPosition_49),
    .io_spriteXPosition_50(graphicEngineVGA_io_spriteXPosition_50),
    .io_spriteXPosition_51(graphicEngineVGA_io_spriteXPosition_51),
    .io_spriteXPosition_122(graphicEngineVGA_io_spriteXPosition_122),
    .io_spriteXPosition_123(graphicEngineVGA_io_spriteXPosition_123),
    .io_spriteXPosition_124(graphicEngineVGA_io_spriteXPosition_124),
    .io_spriteXPosition_125(graphicEngineVGA_io_spriteXPosition_125),
    .io_spriteXPosition_126(graphicEngineVGA_io_spriteXPosition_126),
    .io_spriteXPosition_127(graphicEngineVGA_io_spriteXPosition_127),
    .io_spriteYPosition_0(graphicEngineVGA_io_spriteYPosition_0),
    .io_spriteYPosition_1(graphicEngineVGA_io_spriteYPosition_1),
    .io_spriteYPosition_2(graphicEngineVGA_io_spriteYPosition_2),
    .io_spriteYPosition_3(graphicEngineVGA_io_spriteYPosition_3),
    .io_spriteYPosition_4(graphicEngineVGA_io_spriteYPosition_4),
    .io_spriteYPosition_5(graphicEngineVGA_io_spriteYPosition_5),
    .io_spriteYPosition_6(graphicEngineVGA_io_spriteYPosition_6),
    .io_spriteYPosition_7(graphicEngineVGA_io_spriteYPosition_7),
    .io_spriteYPosition_8(graphicEngineVGA_io_spriteYPosition_8),
    .io_spriteYPosition_9(graphicEngineVGA_io_spriteYPosition_9),
    .io_spriteYPosition_10(graphicEngineVGA_io_spriteYPosition_10),
    .io_spriteYPosition_11(graphicEngineVGA_io_spriteYPosition_11),
    .io_spriteYPosition_12(graphicEngineVGA_io_spriteYPosition_12),
    .io_spriteYPosition_13(graphicEngineVGA_io_spriteYPosition_13),
    .io_spriteYPosition_14(graphicEngineVGA_io_spriteYPosition_14),
    .io_spriteYPosition_15(graphicEngineVGA_io_spriteYPosition_15),
    .io_spriteYPosition_16(graphicEngineVGA_io_spriteYPosition_16),
    .io_spriteYPosition_17(graphicEngineVGA_io_spriteYPosition_17),
    .io_spriteYPosition_18(graphicEngineVGA_io_spriteYPosition_18),
    .io_spriteYPosition_19(graphicEngineVGA_io_spriteYPosition_19),
    .io_spriteYPosition_20(graphicEngineVGA_io_spriteYPosition_20),
    .io_spriteYPosition_21(graphicEngineVGA_io_spriteYPosition_21),
    .io_spriteYPosition_22(graphicEngineVGA_io_spriteYPosition_22),
    .io_spriteYPosition_23(graphicEngineVGA_io_spriteYPosition_23),
    .io_spriteYPosition_24(graphicEngineVGA_io_spriteYPosition_24),
    .io_spriteYPosition_25(graphicEngineVGA_io_spriteYPosition_25),
    .io_spriteYPosition_26(graphicEngineVGA_io_spriteYPosition_26),
    .io_spriteYPosition_27(graphicEngineVGA_io_spriteYPosition_27),
    .io_spriteYPosition_28(graphicEngineVGA_io_spriteYPosition_28),
    .io_spriteYPosition_29(graphicEngineVGA_io_spriteYPosition_29),
    .io_spriteYPosition_30(graphicEngineVGA_io_spriteYPosition_30),
    .io_spriteYPosition_31(graphicEngineVGA_io_spriteYPosition_31),
    .io_spriteYPosition_32(graphicEngineVGA_io_spriteYPosition_32),
    .io_spriteYPosition_33(graphicEngineVGA_io_spriteYPosition_33),
    .io_spriteYPosition_41(graphicEngineVGA_io_spriteYPosition_41),
    .io_spriteYPosition_42(graphicEngineVGA_io_spriteYPosition_42),
    .io_spriteYPosition_43(graphicEngineVGA_io_spriteYPosition_43),
    .io_spriteYPosition_122(graphicEngineVGA_io_spriteYPosition_122),
    .io_spriteYPosition_123(graphicEngineVGA_io_spriteYPosition_123),
    .io_spriteYPosition_124(graphicEngineVGA_io_spriteYPosition_124),
    .io_spriteYPosition_125(graphicEngineVGA_io_spriteYPosition_125),
    .io_spriteYPosition_126(graphicEngineVGA_io_spriteYPosition_126),
    .io_spriteYPosition_127(graphicEngineVGA_io_spriteYPosition_127),
    .io_spriteVisible_0(graphicEngineVGA_io_spriteVisible_0),
    .io_spriteVisible_1(graphicEngineVGA_io_spriteVisible_1),
    .io_spriteVisible_2(graphicEngineVGA_io_spriteVisible_2),
    .io_spriteVisible_3(graphicEngineVGA_io_spriteVisible_3),
    .io_spriteVisible_4(graphicEngineVGA_io_spriteVisible_4),
    .io_spriteVisible_5(graphicEngineVGA_io_spriteVisible_5),
    .io_spriteVisible_6(graphicEngineVGA_io_spriteVisible_6),
    .io_spriteVisible_7(graphicEngineVGA_io_spriteVisible_7),
    .io_spriteVisible_8(graphicEngineVGA_io_spriteVisible_8),
    .io_spriteVisible_9(graphicEngineVGA_io_spriteVisible_9),
    .io_spriteVisible_10(graphicEngineVGA_io_spriteVisible_10),
    .io_spriteVisible_11(graphicEngineVGA_io_spriteVisible_11),
    .io_spriteVisible_12(graphicEngineVGA_io_spriteVisible_12),
    .io_spriteVisible_13(graphicEngineVGA_io_spriteVisible_13),
    .io_spriteVisible_14(graphicEngineVGA_io_spriteVisible_14),
    .io_spriteVisible_15(graphicEngineVGA_io_spriteVisible_15),
    .io_spriteVisible_16(graphicEngineVGA_io_spriteVisible_16),
    .io_spriteVisible_17(graphicEngineVGA_io_spriteVisible_17),
    .io_spriteVisible_18(graphicEngineVGA_io_spriteVisible_18),
    .io_spriteVisible_19(graphicEngineVGA_io_spriteVisible_19),
    .io_spriteVisible_20(graphicEngineVGA_io_spriteVisible_20),
    .io_spriteVisible_21(graphicEngineVGA_io_spriteVisible_21),
    .io_spriteVisible_22(graphicEngineVGA_io_spriteVisible_22),
    .io_spriteVisible_23(graphicEngineVGA_io_spriteVisible_23),
    .io_spriteVisible_24(graphicEngineVGA_io_spriteVisible_24),
    .io_spriteVisible_25(graphicEngineVGA_io_spriteVisible_25),
    .io_spriteVisible_26(graphicEngineVGA_io_spriteVisible_26),
    .io_spriteVisible_27(graphicEngineVGA_io_spriteVisible_27),
    .io_spriteVisible_28(graphicEngineVGA_io_spriteVisible_28),
    .io_spriteVisible_29(graphicEngineVGA_io_spriteVisible_29),
    .io_spriteVisible_30(graphicEngineVGA_io_spriteVisible_30),
    .io_spriteVisible_31(graphicEngineVGA_io_spriteVisible_31),
    .io_spriteVisible_32(graphicEngineVGA_io_spriteVisible_32),
    .io_spriteVisible_33(graphicEngineVGA_io_spriteVisible_33),
    .io_spriteVisible_41(graphicEngineVGA_io_spriteVisible_41),
    .io_spriteVisible_42(graphicEngineVGA_io_spriteVisible_42),
    .io_spriteVisible_43(graphicEngineVGA_io_spriteVisible_43),
    .io_spriteVisible_44(graphicEngineVGA_io_spriteVisible_44),
    .io_spriteVisible_45(graphicEngineVGA_io_spriteVisible_45),
    .io_spriteVisible_46(graphicEngineVGA_io_spriteVisible_46),
    .io_spriteVisible_47(graphicEngineVGA_io_spriteVisible_47),
    .io_spriteVisible_48(graphicEngineVGA_io_spriteVisible_48),
    .io_spriteVisible_49(graphicEngineVGA_io_spriteVisible_49),
    .io_spriteVisible_50(graphicEngineVGA_io_spriteVisible_50),
    .io_spriteVisible_51(graphicEngineVGA_io_spriteVisible_51),
    .io_spriteVisible_55(graphicEngineVGA_io_spriteVisible_55),
    .io_spriteVisible_56(graphicEngineVGA_io_spriteVisible_56),
    .io_spriteVisible_57(graphicEngineVGA_io_spriteVisible_57),
    .io_spriteVisible_61(graphicEngineVGA_io_spriteVisible_61),
    .io_spriteVisible_62(graphicEngineVGA_io_spriteVisible_62),
    .io_spriteVisible_63(graphicEngineVGA_io_spriteVisible_63),
    .io_spriteVisible_64(graphicEngineVGA_io_spriteVisible_64),
    .io_spriteVisible_65(graphicEngineVGA_io_spriteVisible_65),
    .io_spriteVisible_66(graphicEngineVGA_io_spriteVisible_66),
    .io_spriteVisible_70(graphicEngineVGA_io_spriteVisible_70),
    .io_spriteVisible_71(graphicEngineVGA_io_spriteVisible_71),
    .io_spriteVisible_72(graphicEngineVGA_io_spriteVisible_72),
    .io_spriteFlipVertical_122(graphicEngineVGA_io_spriteFlipVertical_122),
    .io_spriteFlipVertical_123(graphicEngineVGA_io_spriteFlipVertical_123),
    .io_spriteFlipVertical_124(graphicEngineVGA_io_spriteFlipVertical_124),
    .io_spriteFlipVertical_125(graphicEngineVGA_io_spriteFlipVertical_125),
    .io_spriteFlipVertical_126(graphicEngineVGA_io_spriteFlipVertical_126),
    .io_spriteFlipVertical_127(graphicEngineVGA_io_spriteFlipVertical_127),
    .io_viewBoxX_0(graphicEngineVGA_io_viewBoxX_0),
    .io_backBufferWriteData(graphicEngineVGA_io_backBufferWriteData),
    .io_backBufferWriteAddress(graphicEngineVGA_io_backBufferWriteAddress),
    .io_backBufferWriteEnable(graphicEngineVGA_io_backBufferWriteEnable),
    .io_newFrame(graphicEngineVGA_io_newFrame),
    .io_frameUpdateDone(graphicEngineVGA_io_frameUpdateDone),
    .io_missingFrameError(graphicEngineVGA_io_missingFrameError),
    .io_backBufferWriteError(graphicEngineVGA_io_backBufferWriteError),
    .io_viewBoxOutOfRangeError(graphicEngineVGA_io_viewBoxOutOfRangeError),
    .io_vgaRed(graphicEngineVGA_io_vgaRed),
    .io_vgaBlue(graphicEngineVGA_io_vgaBlue),
    .io_vgaGreen(graphicEngineVGA_io_vgaGreen),
    .io_Hsync(graphicEngineVGA_io_Hsync),
    .io_Vsync(graphicEngineVGA_io_Vsync)
  );
  SoundEngine soundEngine ( // @[GameTop.scala 48:27]
    .clock(soundEngine_clock),
    .reset(soundEngine_reset),
    .io_output_0(soundEngine_io_output_0),
    .io_input(soundEngine_io_input)
  );
  GameLogic gameLogic ( // @[GameTop.scala 52:25]
    .clock(gameLogic_clock),
    .reset(gameLogic_reset),
    .io_btnC(gameLogic_io_btnC),
    .io_btnU(gameLogic_io_btnU),
    .io_btnL(gameLogic_io_btnL),
    .io_btnR(gameLogic_io_btnR),
    .io_btnD(gameLogic_io_btnD),
    .io_sw_0(gameLogic_io_sw_0),
    .io_sw_1(gameLogic_io_sw_1),
    .io_sw_2(gameLogic_io_sw_2),
    .io_sw_7(gameLogic_io_sw_7),
    .io_songInput(gameLogic_io_songInput),
    .io_spriteXPosition_0(gameLogic_io_spriteXPosition_0),
    .io_spriteXPosition_1(gameLogic_io_spriteXPosition_1),
    .io_spriteXPosition_2(gameLogic_io_spriteXPosition_2),
    .io_spriteXPosition_3(gameLogic_io_spriteXPosition_3),
    .io_spriteXPosition_4(gameLogic_io_spriteXPosition_4),
    .io_spriteXPosition_5(gameLogic_io_spriteXPosition_5),
    .io_spriteXPosition_6(gameLogic_io_spriteXPosition_6),
    .io_spriteXPosition_7(gameLogic_io_spriteXPosition_7),
    .io_spriteXPosition_8(gameLogic_io_spriteXPosition_8),
    .io_spriteXPosition_9(gameLogic_io_spriteXPosition_9),
    .io_spriteXPosition_10(gameLogic_io_spriteXPosition_10),
    .io_spriteXPosition_11(gameLogic_io_spriteXPosition_11),
    .io_spriteXPosition_12(gameLogic_io_spriteXPosition_12),
    .io_spriteXPosition_13(gameLogic_io_spriteXPosition_13),
    .io_spriteXPosition_14(gameLogic_io_spriteXPosition_14),
    .io_spriteXPosition_15(gameLogic_io_spriteXPosition_15),
    .io_spriteXPosition_16(gameLogic_io_spriteXPosition_16),
    .io_spriteXPosition_17(gameLogic_io_spriteXPosition_17),
    .io_spriteXPosition_18(gameLogic_io_spriteXPosition_18),
    .io_spriteXPosition_19(gameLogic_io_spriteXPosition_19),
    .io_spriteXPosition_20(gameLogic_io_spriteXPosition_20),
    .io_spriteXPosition_21(gameLogic_io_spriteXPosition_21),
    .io_spriteXPosition_22(gameLogic_io_spriteXPosition_22),
    .io_spriteXPosition_23(gameLogic_io_spriteXPosition_23),
    .io_spriteXPosition_24(gameLogic_io_spriteXPosition_24),
    .io_spriteXPosition_25(gameLogic_io_spriteXPosition_25),
    .io_spriteXPosition_26(gameLogic_io_spriteXPosition_26),
    .io_spriteXPosition_27(gameLogic_io_spriteXPosition_27),
    .io_spriteXPosition_28(gameLogic_io_spriteXPosition_28),
    .io_spriteXPosition_29(gameLogic_io_spriteXPosition_29),
    .io_spriteXPosition_30(gameLogic_io_spriteXPosition_30),
    .io_spriteXPosition_31(gameLogic_io_spriteXPosition_31),
    .io_spriteXPosition_32(gameLogic_io_spriteXPosition_32),
    .io_spriteXPosition_33(gameLogic_io_spriteXPosition_33),
    .io_spriteXPosition_41(gameLogic_io_spriteXPosition_41),
    .io_spriteXPosition_42(gameLogic_io_spriteXPosition_42),
    .io_spriteXPosition_43(gameLogic_io_spriteXPosition_43),
    .io_spriteXPosition_44(gameLogic_io_spriteXPosition_44),
    .io_spriteXPosition_45(gameLogic_io_spriteXPosition_45),
    .io_spriteXPosition_46(gameLogic_io_spriteXPosition_46),
    .io_spriteXPosition_47(gameLogic_io_spriteXPosition_47),
    .io_spriteXPosition_48(gameLogic_io_spriteXPosition_48),
    .io_spriteXPosition_49(gameLogic_io_spriteXPosition_49),
    .io_spriteXPosition_50(gameLogic_io_spriteXPosition_50),
    .io_spriteXPosition_51(gameLogic_io_spriteXPosition_51),
    .io_spriteXPosition_122(gameLogic_io_spriteXPosition_122),
    .io_spriteXPosition_123(gameLogic_io_spriteXPosition_123),
    .io_spriteXPosition_124(gameLogic_io_spriteXPosition_124),
    .io_spriteXPosition_125(gameLogic_io_spriteXPosition_125),
    .io_spriteXPosition_126(gameLogic_io_spriteXPosition_126),
    .io_spriteXPosition_127(gameLogic_io_spriteXPosition_127),
    .io_spriteYPosition_0(gameLogic_io_spriteYPosition_0),
    .io_spriteYPosition_1(gameLogic_io_spriteYPosition_1),
    .io_spriteYPosition_2(gameLogic_io_spriteYPosition_2),
    .io_spriteYPosition_3(gameLogic_io_spriteYPosition_3),
    .io_spriteYPosition_4(gameLogic_io_spriteYPosition_4),
    .io_spriteYPosition_5(gameLogic_io_spriteYPosition_5),
    .io_spriteYPosition_6(gameLogic_io_spriteYPosition_6),
    .io_spriteYPosition_7(gameLogic_io_spriteYPosition_7),
    .io_spriteYPosition_8(gameLogic_io_spriteYPosition_8),
    .io_spriteYPosition_9(gameLogic_io_spriteYPosition_9),
    .io_spriteYPosition_10(gameLogic_io_spriteYPosition_10),
    .io_spriteYPosition_11(gameLogic_io_spriteYPosition_11),
    .io_spriteYPosition_12(gameLogic_io_spriteYPosition_12),
    .io_spriteYPosition_13(gameLogic_io_spriteYPosition_13),
    .io_spriteYPosition_14(gameLogic_io_spriteYPosition_14),
    .io_spriteYPosition_15(gameLogic_io_spriteYPosition_15),
    .io_spriteYPosition_16(gameLogic_io_spriteYPosition_16),
    .io_spriteYPosition_17(gameLogic_io_spriteYPosition_17),
    .io_spriteYPosition_18(gameLogic_io_spriteYPosition_18),
    .io_spriteYPosition_19(gameLogic_io_spriteYPosition_19),
    .io_spriteYPosition_20(gameLogic_io_spriteYPosition_20),
    .io_spriteYPosition_21(gameLogic_io_spriteYPosition_21),
    .io_spriteYPosition_22(gameLogic_io_spriteYPosition_22),
    .io_spriteYPosition_23(gameLogic_io_spriteYPosition_23),
    .io_spriteYPosition_24(gameLogic_io_spriteYPosition_24),
    .io_spriteYPosition_25(gameLogic_io_spriteYPosition_25),
    .io_spriteYPosition_26(gameLogic_io_spriteYPosition_26),
    .io_spriteYPosition_27(gameLogic_io_spriteYPosition_27),
    .io_spriteYPosition_28(gameLogic_io_spriteYPosition_28),
    .io_spriteYPosition_29(gameLogic_io_spriteYPosition_29),
    .io_spriteYPosition_30(gameLogic_io_spriteYPosition_30),
    .io_spriteYPosition_31(gameLogic_io_spriteYPosition_31),
    .io_spriteYPosition_32(gameLogic_io_spriteYPosition_32),
    .io_spriteYPosition_33(gameLogic_io_spriteYPosition_33),
    .io_spriteYPosition_41(gameLogic_io_spriteYPosition_41),
    .io_spriteYPosition_42(gameLogic_io_spriteYPosition_42),
    .io_spriteYPosition_43(gameLogic_io_spriteYPosition_43),
    .io_spriteYPosition_122(gameLogic_io_spriteYPosition_122),
    .io_spriteYPosition_123(gameLogic_io_spriteYPosition_123),
    .io_spriteYPosition_124(gameLogic_io_spriteYPosition_124),
    .io_spriteYPosition_125(gameLogic_io_spriteYPosition_125),
    .io_spriteYPosition_126(gameLogic_io_spriteYPosition_126),
    .io_spriteYPosition_127(gameLogic_io_spriteYPosition_127),
    .io_spriteVisible_0(gameLogic_io_spriteVisible_0),
    .io_spriteVisible_1(gameLogic_io_spriteVisible_1),
    .io_spriteVisible_2(gameLogic_io_spriteVisible_2),
    .io_spriteVisible_3(gameLogic_io_spriteVisible_3),
    .io_spriteVisible_4(gameLogic_io_spriteVisible_4),
    .io_spriteVisible_5(gameLogic_io_spriteVisible_5),
    .io_spriteVisible_6(gameLogic_io_spriteVisible_6),
    .io_spriteVisible_7(gameLogic_io_spriteVisible_7),
    .io_spriteVisible_8(gameLogic_io_spriteVisible_8),
    .io_spriteVisible_9(gameLogic_io_spriteVisible_9),
    .io_spriteVisible_10(gameLogic_io_spriteVisible_10),
    .io_spriteVisible_11(gameLogic_io_spriteVisible_11),
    .io_spriteVisible_12(gameLogic_io_spriteVisible_12),
    .io_spriteVisible_13(gameLogic_io_spriteVisible_13),
    .io_spriteVisible_14(gameLogic_io_spriteVisible_14),
    .io_spriteVisible_15(gameLogic_io_spriteVisible_15),
    .io_spriteVisible_16(gameLogic_io_spriteVisible_16),
    .io_spriteVisible_17(gameLogic_io_spriteVisible_17),
    .io_spriteVisible_18(gameLogic_io_spriteVisible_18),
    .io_spriteVisible_19(gameLogic_io_spriteVisible_19),
    .io_spriteVisible_20(gameLogic_io_spriteVisible_20),
    .io_spriteVisible_21(gameLogic_io_spriteVisible_21),
    .io_spriteVisible_22(gameLogic_io_spriteVisible_22),
    .io_spriteVisible_23(gameLogic_io_spriteVisible_23),
    .io_spriteVisible_24(gameLogic_io_spriteVisible_24),
    .io_spriteVisible_25(gameLogic_io_spriteVisible_25),
    .io_spriteVisible_26(gameLogic_io_spriteVisible_26),
    .io_spriteVisible_27(gameLogic_io_spriteVisible_27),
    .io_spriteVisible_28(gameLogic_io_spriteVisible_28),
    .io_spriteVisible_29(gameLogic_io_spriteVisible_29),
    .io_spriteVisible_30(gameLogic_io_spriteVisible_30),
    .io_spriteVisible_31(gameLogic_io_spriteVisible_31),
    .io_spriteVisible_32(gameLogic_io_spriteVisible_32),
    .io_spriteVisible_33(gameLogic_io_spriteVisible_33),
    .io_spriteVisible_41(gameLogic_io_spriteVisible_41),
    .io_spriteVisible_42(gameLogic_io_spriteVisible_42),
    .io_spriteVisible_43(gameLogic_io_spriteVisible_43),
    .io_spriteVisible_44(gameLogic_io_spriteVisible_44),
    .io_spriteVisible_45(gameLogic_io_spriteVisible_45),
    .io_spriteVisible_46(gameLogic_io_spriteVisible_46),
    .io_spriteVisible_47(gameLogic_io_spriteVisible_47),
    .io_spriteVisible_48(gameLogic_io_spriteVisible_48),
    .io_spriteVisible_49(gameLogic_io_spriteVisible_49),
    .io_spriteVisible_50(gameLogic_io_spriteVisible_50),
    .io_spriteVisible_51(gameLogic_io_spriteVisible_51),
    .io_spriteVisible_55(gameLogic_io_spriteVisible_55),
    .io_spriteVisible_56(gameLogic_io_spriteVisible_56),
    .io_spriteVisible_57(gameLogic_io_spriteVisible_57),
    .io_spriteVisible_61(gameLogic_io_spriteVisible_61),
    .io_spriteVisible_62(gameLogic_io_spriteVisible_62),
    .io_spriteVisible_63(gameLogic_io_spriteVisible_63),
    .io_spriteVisible_64(gameLogic_io_spriteVisible_64),
    .io_spriteVisible_65(gameLogic_io_spriteVisible_65),
    .io_spriteVisible_66(gameLogic_io_spriteVisible_66),
    .io_spriteVisible_70(gameLogic_io_spriteVisible_70),
    .io_spriteVisible_71(gameLogic_io_spriteVisible_71),
    .io_spriteVisible_72(gameLogic_io_spriteVisible_72),
    .io_spriteFlipVertical_122(gameLogic_io_spriteFlipVertical_122),
    .io_spriteFlipVertical_123(gameLogic_io_spriteFlipVertical_123),
    .io_spriteFlipVertical_124(gameLogic_io_spriteFlipVertical_124),
    .io_spriteFlipVertical_125(gameLogic_io_spriteFlipVertical_125),
    .io_spriteFlipVertical_126(gameLogic_io_spriteFlipVertical_126),
    .io_spriteFlipVertical_127(gameLogic_io_spriteFlipVertical_127),
    .io_viewBoxX_0(gameLogic_io_viewBoxX_0),
    .io_backBufferWriteData(gameLogic_io_backBufferWriteData),
    .io_backBufferWriteAddress(gameLogic_io_backBufferWriteAddress),
    .io_backBufferWriteEnable(gameLogic_io_backBufferWriteEnable),
    .io_newFrame(gameLogic_io_newFrame),
    .io_frameUpdateDone(gameLogic_io_frameUpdateDone)
  );
  assign io_vgaRed = graphicEngineVGA_io_vgaRed; // @[GameTop.scala 110:13]
  assign io_vgaBlue = graphicEngineVGA_io_vgaBlue; // @[GameTop.scala 112:14]
  assign io_vgaGreen = graphicEngineVGA_io_vgaGreen; // @[GameTop.scala 111:15]
  assign io_Hsync = graphicEngineVGA_io_Hsync; // @[GameTop.scala 113:12]
  assign io_Vsync = graphicEngineVGA_io_Vsync; // @[GameTop.scala 114:12]
  assign io_soundOutput_0 = soundEngine_io_output_0; // @[GameTop.scala 68:18]
  assign io_missingFrameError = graphicEngineVGA_io_missingFrameError; // @[GameTop.scala 125:24]
  assign io_backBufferWriteError = graphicEngineVGA_io_backBufferWriteError; // @[GameTop.scala 126:27]
  assign io_viewBoxOutOfRangeError = graphicEngineVGA_io_viewBoxOutOfRangeError; // @[GameTop.scala 127:29]
  assign graphicEngineVGA_clock = clock;
  assign graphicEngineVGA_reset = _T_3 ? 1'h0 : 1'h1; // @[GameTop.scala 94:26]
  assign graphicEngineVGA_io_spriteXPosition_0 = gameLogic_io_spriteXPosition_0; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_1 = gameLogic_io_spriteXPosition_1; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_2 = gameLogic_io_spriteXPosition_2; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_3 = gameLogic_io_spriteXPosition_3; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_4 = gameLogic_io_spriteXPosition_4; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_5 = gameLogic_io_spriteXPosition_5; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_6 = gameLogic_io_spriteXPosition_6; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_7 = gameLogic_io_spriteXPosition_7; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_8 = gameLogic_io_spriteXPosition_8; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_9 = gameLogic_io_spriteXPosition_9; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_10 = gameLogic_io_spriteXPosition_10; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_11 = gameLogic_io_spriteXPosition_11; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_12 = gameLogic_io_spriteXPosition_12; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_13 = gameLogic_io_spriteXPosition_13; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_14 = gameLogic_io_spriteXPosition_14; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_15 = gameLogic_io_spriteXPosition_15; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_16 = gameLogic_io_spriteXPosition_16; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_17 = gameLogic_io_spriteXPosition_17; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_18 = gameLogic_io_spriteXPosition_18; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_19 = gameLogic_io_spriteXPosition_19; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_20 = gameLogic_io_spriteXPosition_20; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_21 = gameLogic_io_spriteXPosition_21; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_22 = gameLogic_io_spriteXPosition_22; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_23 = gameLogic_io_spriteXPosition_23; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_24 = gameLogic_io_spriteXPosition_24; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_25 = gameLogic_io_spriteXPosition_25; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_26 = gameLogic_io_spriteXPosition_26; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_27 = gameLogic_io_spriteXPosition_27; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_28 = gameLogic_io_spriteXPosition_28; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_29 = gameLogic_io_spriteXPosition_29; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_30 = gameLogic_io_spriteXPosition_30; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_31 = gameLogic_io_spriteXPosition_31; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_32 = gameLogic_io_spriteXPosition_32; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_33 = gameLogic_io_spriteXPosition_33; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_41 = gameLogic_io_spriteXPosition_41; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_42 = gameLogic_io_spriteXPosition_42; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_43 = gameLogic_io_spriteXPosition_43; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_44 = gameLogic_io_spriteXPosition_44; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_45 = gameLogic_io_spriteXPosition_45; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_46 = gameLogic_io_spriteXPosition_46; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_47 = gameLogic_io_spriteXPosition_47; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_48 = gameLogic_io_spriteXPosition_48; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_49 = gameLogic_io_spriteXPosition_49; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_50 = gameLogic_io_spriteXPosition_50; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_51 = gameLogic_io_spriteXPosition_51; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_122 = gameLogic_io_spriteXPosition_122; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_123 = gameLogic_io_spriteXPosition_123; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_124 = gameLogic_io_spriteXPosition_124; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_125 = gameLogic_io_spriteXPosition_125; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_126 = gameLogic_io_spriteXPosition_126; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteXPosition_127 = gameLogic_io_spriteXPosition_127; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_0 = gameLogic_io_spriteYPosition_0; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_1 = gameLogic_io_spriteYPosition_1; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_2 = gameLogic_io_spriteYPosition_2; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_3 = gameLogic_io_spriteYPosition_3; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_4 = gameLogic_io_spriteYPosition_4; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_5 = gameLogic_io_spriteYPosition_5; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_6 = gameLogic_io_spriteYPosition_6; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_7 = gameLogic_io_spriteYPosition_7; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_8 = gameLogic_io_spriteYPosition_8; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_9 = gameLogic_io_spriteYPosition_9; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_10 = gameLogic_io_spriteYPosition_10; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_11 = gameLogic_io_spriteYPosition_11; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_12 = gameLogic_io_spriteYPosition_12; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_13 = gameLogic_io_spriteYPosition_13; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_14 = gameLogic_io_spriteYPosition_14; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_15 = gameLogic_io_spriteYPosition_15; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_16 = gameLogic_io_spriteYPosition_16; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_17 = gameLogic_io_spriteYPosition_17; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_18 = gameLogic_io_spriteYPosition_18; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_19 = gameLogic_io_spriteYPosition_19; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_20 = gameLogic_io_spriteYPosition_20; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_21 = gameLogic_io_spriteYPosition_21; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_22 = gameLogic_io_spriteYPosition_22; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_23 = gameLogic_io_spriteYPosition_23; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_24 = gameLogic_io_spriteYPosition_24; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_25 = gameLogic_io_spriteYPosition_25; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_26 = gameLogic_io_spriteYPosition_26; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_27 = gameLogic_io_spriteYPosition_27; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_28 = gameLogic_io_spriteYPosition_28; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_29 = gameLogic_io_spriteYPosition_29; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_30 = gameLogic_io_spriteYPosition_30; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_31 = gameLogic_io_spriteYPosition_31; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_32 = gameLogic_io_spriteYPosition_32; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_33 = gameLogic_io_spriteYPosition_33; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_41 = gameLogic_io_spriteYPosition_41; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_42 = gameLogic_io_spriteYPosition_42; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_43 = gameLogic_io_spriteYPosition_43; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_122 = gameLogic_io_spriteYPosition_122; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_123 = gameLogic_io_spriteYPosition_123; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_124 = gameLogic_io_spriteYPosition_124; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_125 = gameLogic_io_spriteYPosition_125; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_126 = gameLogic_io_spriteYPosition_126; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteYPosition_127 = gameLogic_io_spriteYPosition_127; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteVisible_0 = gameLogic_io_spriteVisible_0; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_1 = gameLogic_io_spriteVisible_1; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_2 = gameLogic_io_spriteVisible_2; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_3 = gameLogic_io_spriteVisible_3; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_4 = gameLogic_io_spriteVisible_4; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_5 = gameLogic_io_spriteVisible_5; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_6 = gameLogic_io_spriteVisible_6; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_7 = gameLogic_io_spriteVisible_7; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_8 = gameLogic_io_spriteVisible_8; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_9 = gameLogic_io_spriteVisible_9; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_10 = gameLogic_io_spriteVisible_10; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_11 = gameLogic_io_spriteVisible_11; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_12 = gameLogic_io_spriteVisible_12; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_13 = gameLogic_io_spriteVisible_13; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_14 = gameLogic_io_spriteVisible_14; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_15 = gameLogic_io_spriteVisible_15; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_16 = gameLogic_io_spriteVisible_16; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_17 = gameLogic_io_spriteVisible_17; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_18 = gameLogic_io_spriteVisible_18; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_19 = gameLogic_io_spriteVisible_19; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_20 = gameLogic_io_spriteVisible_20; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_21 = gameLogic_io_spriteVisible_21; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_22 = gameLogic_io_spriteVisible_22; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_23 = gameLogic_io_spriteVisible_23; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_24 = gameLogic_io_spriteVisible_24; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_25 = gameLogic_io_spriteVisible_25; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_26 = gameLogic_io_spriteVisible_26; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_27 = gameLogic_io_spriteVisible_27; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_28 = gameLogic_io_spriteVisible_28; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_29 = gameLogic_io_spriteVisible_29; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_30 = gameLogic_io_spriteVisible_30; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_31 = gameLogic_io_spriteVisible_31; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_32 = gameLogic_io_spriteVisible_32; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_33 = gameLogic_io_spriteVisible_33; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_41 = gameLogic_io_spriteVisible_41; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_42 = gameLogic_io_spriteVisible_42; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_43 = gameLogic_io_spriteVisible_43; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_44 = gameLogic_io_spriteVisible_44; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_45 = gameLogic_io_spriteVisible_45; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_46 = gameLogic_io_spriteVisible_46; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_47 = gameLogic_io_spriteVisible_47; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_48 = gameLogic_io_spriteVisible_48; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_49 = gameLogic_io_spriteVisible_49; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_50 = gameLogic_io_spriteVisible_50; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_51 = gameLogic_io_spriteVisible_51; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_55 = gameLogic_io_spriteVisible_55; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_56 = gameLogic_io_spriteVisible_56; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_57 = gameLogic_io_spriteVisible_57; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_61 = gameLogic_io_spriteVisible_61; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_62 = gameLogic_io_spriteVisible_62; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_63 = gameLogic_io_spriteVisible_63; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_64 = gameLogic_io_spriteVisible_64; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_65 = gameLogic_io_spriteVisible_65; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_66 = gameLogic_io_spriteVisible_66; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_70 = gameLogic_io_spriteVisible_70; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_71 = gameLogic_io_spriteVisible_71; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteVisible_72 = gameLogic_io_spriteVisible_72; // @[GameTop.scala 132:37]
  assign graphicEngineVGA_io_spriteFlipVertical_122 = gameLogic_io_spriteFlipVertical_122; // @[GameTop.scala 135:42]
  assign graphicEngineVGA_io_spriteFlipVertical_123 = gameLogic_io_spriteFlipVertical_123; // @[GameTop.scala 135:42]
  assign graphicEngineVGA_io_spriteFlipVertical_124 = gameLogic_io_spriteFlipVertical_124; // @[GameTop.scala 135:42]
  assign graphicEngineVGA_io_spriteFlipVertical_125 = gameLogic_io_spriteFlipVertical_125; // @[GameTop.scala 135:42]
  assign graphicEngineVGA_io_spriteFlipVertical_126 = gameLogic_io_spriteFlipVertical_126; // @[GameTop.scala 135:42]
  assign graphicEngineVGA_io_spriteFlipVertical_127 = gameLogic_io_spriteFlipVertical_127; // @[GameTop.scala 135:42]
  assign graphicEngineVGA_io_viewBoxX_0 = gameLogic_io_viewBoxX_0; // @[GameTop.scala 144:32]
  assign graphicEngineVGA_io_backBufferWriteData = gameLogic_io_backBufferWriteData; // @[GameTop.scala 148:43]
  assign graphicEngineVGA_io_backBufferWriteAddress = gameLogic_io_backBufferWriteAddress; // @[GameTop.scala 149:46]
  assign graphicEngineVGA_io_backBufferWriteEnable = gameLogic_io_backBufferWriteEnable; // @[GameTop.scala 150:45]
  assign graphicEngineVGA_io_frameUpdateDone = gameLogic_io_frameUpdateDone; // @[GameTop.scala 154:39]
  assign soundEngine_clock = clock;
  assign soundEngine_reset = reset;
  assign soundEngine_io_input = gameLogic_io_songInput; // @[GameTop.scala 65:24]
  assign gameLogic_clock = clock;
  assign gameLogic_reset = _T_3 ? 1'h0 : 1'h1; // @[GameTop.scala 95:19]
  assign gameLogic_io_btnC = btnCState; // @[GameTop.scala 103:21]
  assign gameLogic_io_btnU = btnUState; // @[GameTop.scala 104:21]
  assign gameLogic_io_btnL = btnLState; // @[GameTop.scala 105:21]
  assign gameLogic_io_btnR = btnRState; // @[GameTop.scala 106:21]
  assign gameLogic_io_btnD = btnDState; // @[GameTop.scala 107:21]
  assign gameLogic_io_sw_0 = _T_18; // @[GameTop.scala 118:24]
  assign gameLogic_io_sw_1 = _T_21; // @[GameTop.scala 118:24]
  assign gameLogic_io_sw_2 = _T_24; // @[GameTop.scala 118:24]
  assign gameLogic_io_sw_7 = _T_39; // @[GameTop.scala 118:24]
  assign gameLogic_io_newFrame = graphicEngineVGA_io_newFrame; // @[GameTop.scala 153:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounceCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  resetReleaseCounter = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  _T_7_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_7_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_7_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btnCState = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_9_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_9_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_9_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btnUState = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_11_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_11_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_11_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btnLState = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_13_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_13_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_13_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btnRState = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_15_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_15_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_15_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  btnDState = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_17_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_17_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_17_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_18 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_20_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_20_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_20_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_21 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_23_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_23_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_23_2 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_24 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_38_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_38_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_38_2 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_39 = _RAND_37[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      debounceCounter <= 21'h0;
    end else if (debounceSampleEn) begin
      debounceCounter <= 21'h0;
    end else begin
      debounceCounter <= _T_2;
    end
    if (reset) begin
      resetReleaseCounter <= 22'h0;
    end else if (!(_T_3)) begin
      resetReleaseCounter <= _T_5;
    end
    if (reset) begin
      _T_7_0 <= 1'h0;
    end else begin
      _T_7_0 <= _T_7_1;
    end
    if (reset) begin
      _T_7_1 <= 1'h0;
    end else begin
      _T_7_1 <= _T_7_2;
    end
    if (reset) begin
      _T_7_2 <= 1'h0;
    end else begin
      _T_7_2 <= io_btnC;
    end
    if (reset) begin
      btnCState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnCState <= _T_7_0;
    end
    if (reset) begin
      _T_9_0 <= 1'h0;
    end else begin
      _T_9_0 <= _T_9_1;
    end
    if (reset) begin
      _T_9_1 <= 1'h0;
    end else begin
      _T_9_1 <= _T_9_2;
    end
    if (reset) begin
      _T_9_2 <= 1'h0;
    end else begin
      _T_9_2 <= io_btnU;
    end
    if (reset) begin
      btnUState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnUState <= _T_9_0;
    end
    if (reset) begin
      _T_11_0 <= 1'h0;
    end else begin
      _T_11_0 <= _T_11_1;
    end
    if (reset) begin
      _T_11_1 <= 1'h0;
    end else begin
      _T_11_1 <= _T_11_2;
    end
    if (reset) begin
      _T_11_2 <= 1'h0;
    end else begin
      _T_11_2 <= io_btnL;
    end
    if (reset) begin
      btnLState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnLState <= _T_11_0;
    end
    if (reset) begin
      _T_13_0 <= 1'h0;
    end else begin
      _T_13_0 <= _T_13_1;
    end
    if (reset) begin
      _T_13_1 <= 1'h0;
    end else begin
      _T_13_1 <= _T_13_2;
    end
    if (reset) begin
      _T_13_2 <= 1'h0;
    end else begin
      _T_13_2 <= io_btnR;
    end
    if (reset) begin
      btnRState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnRState <= _T_13_0;
    end
    if (reset) begin
      _T_15_0 <= 1'h0;
    end else begin
      _T_15_0 <= _T_15_1;
    end
    if (reset) begin
      _T_15_1 <= 1'h0;
    end else begin
      _T_15_1 <= _T_15_2;
    end
    if (reset) begin
      _T_15_2 <= 1'h0;
    end else begin
      _T_15_2 <= io_btnD;
    end
    if (reset) begin
      btnDState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnDState <= _T_15_0;
    end
    if (reset) begin
      _T_17_0 <= 1'h0;
    end else begin
      _T_17_0 <= _T_17_1;
    end
    if (reset) begin
      _T_17_1 <= 1'h0;
    end else begin
      _T_17_1 <= _T_17_2;
    end
    if (reset) begin
      _T_17_2 <= 1'h0;
    end else begin
      _T_17_2 <= io_sw_0;
    end
    if (reset) begin
      _T_18 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_18 <= _T_17_0;
    end
    if (reset) begin
      _T_20_0 <= 1'h0;
    end else begin
      _T_20_0 <= _T_20_1;
    end
    if (reset) begin
      _T_20_1 <= 1'h0;
    end else begin
      _T_20_1 <= _T_20_2;
    end
    if (reset) begin
      _T_20_2 <= 1'h0;
    end else begin
      _T_20_2 <= io_sw_1;
    end
    if (reset) begin
      _T_21 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_21 <= _T_20_0;
    end
    if (reset) begin
      _T_23_0 <= 1'h0;
    end else begin
      _T_23_0 <= _T_23_1;
    end
    if (reset) begin
      _T_23_1 <= 1'h0;
    end else begin
      _T_23_1 <= _T_23_2;
    end
    if (reset) begin
      _T_23_2 <= 1'h0;
    end else begin
      _T_23_2 <= io_sw_2;
    end
    if (reset) begin
      _T_24 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_24 <= _T_23_0;
    end
    if (reset) begin
      _T_38_0 <= 1'h0;
    end else begin
      _T_38_0 <= _T_38_1;
    end
    if (reset) begin
      _T_38_1 <= 1'h0;
    end else begin
      _T_38_1 <= _T_38_2;
    end
    if (reset) begin
      _T_38_2 <= 1'h0;
    end else begin
      _T_38_2 <= io_sw_7;
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_39 <= _T_38_0;
    end
  end
endmodule
module Top(
  input        clock,
  input        reset,
  input        io_btnC,
  input        io_btnU,
  input        io_btnL,
  input        io_btnR,
  input        io_btnD,
  output [3:0] io_vgaRed,
  output [3:0] io_vgaGreen,
  output [3:0] io_vgaBlue,
  output       io_Hsync,
  output       io_Vsync,
  input        io_sw_0,
  input        io_sw_1,
  input        io_sw_2,
  input        io_sw_3,
  input        io_sw_4,
  input        io_sw_5,
  input        io_sw_6,
  input        io_sw_7,
  output       io_led_0,
  output       io_led_1,
  output       io_led_2,
  output       io_led_3,
  output       io_led_4,
  output       io_led_5,
  output       io_led_6,
  output       io_led_7,
  output       io_soundOutput_0,
  output       io_missingFrameError,
  output       io_backBufferWriteError,
  output       io_viewBoxOutOfRangeError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  gameTop_clock; // @[Top.scala 42:23]
  wire  gameTop_reset; // @[Top.scala 42:23]
  wire  gameTop_io_btnC; // @[Top.scala 42:23]
  wire  gameTop_io_btnU; // @[Top.scala 42:23]
  wire  gameTop_io_btnL; // @[Top.scala 42:23]
  wire  gameTop_io_btnR; // @[Top.scala 42:23]
  wire  gameTop_io_btnD; // @[Top.scala 42:23]
  wire [3:0] gameTop_io_vgaRed; // @[Top.scala 42:23]
  wire [3:0] gameTop_io_vgaBlue; // @[Top.scala 42:23]
  wire [3:0] gameTop_io_vgaGreen; // @[Top.scala 42:23]
  wire  gameTop_io_Hsync; // @[Top.scala 42:23]
  wire  gameTop_io_Vsync; // @[Top.scala 42:23]
  wire  gameTop_io_sw_0; // @[Top.scala 42:23]
  wire  gameTop_io_sw_1; // @[Top.scala 42:23]
  wire  gameTop_io_sw_2; // @[Top.scala 42:23]
  wire  gameTop_io_sw_7; // @[Top.scala 42:23]
  wire  gameTop_io_soundOutput_0; // @[Top.scala 42:23]
  wire  gameTop_io_missingFrameError; // @[Top.scala 42:23]
  wire  gameTop_io_backBufferWriteError; // @[Top.scala 42:23]
  wire  gameTop_io_viewBoxOutOfRangeError; // @[Top.scala 42:23]
  reg  _T_1; // @[Top.scala 47:48]
  reg  _T_2; // @[Top.scala 47:40]
  reg  _T_3; // @[Top.scala 47:32]
  reg  pipeResetReg_0; // @[Top.scala 52:25]
  reg  pipeResetReg_1; // @[Top.scala 52:25]
  reg  pipeResetReg_2; // @[Top.scala 52:25]
  reg  pipeResetReg_3; // @[Top.scala 52:25]
  reg  pipeResetReg_4; // @[Top.scala 52:25]
  wire [4:0] _T_7 = {pipeResetReg_4,pipeResetReg_3,pipeResetReg_2,pipeResetReg_1,pipeResetReg_0}; // @[Top.scala 57:33]
  GameTop gameTop ( // @[Top.scala 42:23]
    .clock(gameTop_clock),
    .reset(gameTop_reset),
    .io_btnC(gameTop_io_btnC),
    .io_btnU(gameTop_io_btnU),
    .io_btnL(gameTop_io_btnL),
    .io_btnR(gameTop_io_btnR),
    .io_btnD(gameTop_io_btnD),
    .io_vgaRed(gameTop_io_vgaRed),
    .io_vgaBlue(gameTop_io_vgaBlue),
    .io_vgaGreen(gameTop_io_vgaGreen),
    .io_Hsync(gameTop_io_Hsync),
    .io_Vsync(gameTop_io_Vsync),
    .io_sw_0(gameTop_io_sw_0),
    .io_sw_1(gameTop_io_sw_1),
    .io_sw_2(gameTop_io_sw_2),
    .io_sw_7(gameTop_io_sw_7),
    .io_soundOutput_0(gameTop_io_soundOutput_0),
    .io_missingFrameError(gameTop_io_missingFrameError),
    .io_backBufferWriteError(gameTop_io_backBufferWriteError),
    .io_viewBoxOutOfRangeError(gameTop_io_viewBoxOutOfRangeError)
  );
  assign io_vgaRed = gameTop_io_vgaRed; // @[Top.scala 60:14]
  assign io_vgaGreen = gameTop_io_vgaGreen; // @[Top.scala 60:14]
  assign io_vgaBlue = gameTop_io_vgaBlue; // @[Top.scala 60:14]
  assign io_Hsync = gameTop_io_Hsync; // @[Top.scala 60:14]
  assign io_Vsync = gameTop_io_Vsync; // @[Top.scala 60:14]
  assign io_led_0 = 1'h0; // @[Top.scala 60:14]
  assign io_led_1 = 1'h0; // @[Top.scala 60:14]
  assign io_led_2 = 1'h0; // @[Top.scala 60:14]
  assign io_led_3 = 1'h0; // @[Top.scala 60:14]
  assign io_led_4 = 1'h0; // @[Top.scala 60:14]
  assign io_led_5 = 1'h0; // @[Top.scala 60:14]
  assign io_led_6 = 1'h0; // @[Top.scala 60:14]
  assign io_led_7 = 1'h0; // @[Top.scala 60:14]
  assign io_soundOutput_0 = gameTop_io_soundOutput_0; // @[Top.scala 60:14]
  assign io_missingFrameError = gameTop_io_missingFrameError; // @[Top.scala 60:14]
  assign io_backBufferWriteError = gameTop_io_backBufferWriteError; // @[Top.scala 60:14]
  assign io_viewBoxOutOfRangeError = gameTop_io_viewBoxOutOfRangeError; // @[Top.scala 60:14]
  assign gameTop_clock = clock;
  assign gameTop_reset = |_T_7; // @[Top.scala 57:17]
  assign gameTop_io_btnC = io_btnC; // @[Top.scala 60:14]
  assign gameTop_io_btnU = io_btnU; // @[Top.scala 60:14]
  assign gameTop_io_btnL = io_btnL; // @[Top.scala 60:14]
  assign gameTop_io_btnR = io_btnR; // @[Top.scala 60:14]
  assign gameTop_io_btnD = io_btnD; // @[Top.scala 60:14]
  assign gameTop_io_sw_0 = io_sw_0; // @[Top.scala 60:14]
  assign gameTop_io_sw_1 = io_sw_1; // @[Top.scala 60:14]
  assign gameTop_io_sw_2 = io_sw_2; // @[Top.scala 60:14]
  assign gameTop_io_sw_7 = io_sw_7; // @[Top.scala 60:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_2 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipeResetReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipeResetReg_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pipeResetReg_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipeResetReg_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pipeResetReg_4 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= reset;
    _T_2 <= _T_1;
    _T_3 <= _T_2;
    pipeResetReg_0 <= pipeResetReg_1;
    pipeResetReg_1 <= pipeResetReg_2;
    pipeResetReg_2 <= pipeResetReg_3;
    pipeResetReg_3 <= pipeResetReg_4;
    pipeResetReg_4 <= ~_T_3;
  end
endmodule
