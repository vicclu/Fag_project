module Memory(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_1(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_2(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_3(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_4(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_5(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_6(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_7(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_8(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_8.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_9(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_9.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_10(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_10.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_11(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_11.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_12(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_12.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_13(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_13.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_14(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_14.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_15(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_15.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_16(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_16.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_17(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_17.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_18(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_18.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_19(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_19.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_20(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_20.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_21(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_21.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_22(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_22.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_23(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_23.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_24(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_24.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_25(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_25.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_26(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_26.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_27(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_27.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_28(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_28.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_29(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_29.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_30(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_30.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_31(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_31.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_32(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead,
  input         io_writeEnable,
  input  [4:0]  io_dataWrite
);
  wire  RamSpWf_clk; // @[Memory.scala 57:26]
  wire  RamSpWf_we; // @[Memory.scala 57:26]
  wire  RamSpWf_en; // @[Memory.scala 57:26]
  wire [10:0] RamSpWf_addr; // @[Memory.scala 57:26]
  wire [4:0] RamSpWf_di; // @[Memory.scala 57:26]
  wire [4:0] RamSpWf_dout; // @[Memory.scala 57:26]
  RamSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5)) RamSpWf ( // @[Memory.scala 57:26]
    .clk(RamSpWf_clk),
    .we(RamSpWf_we),
    .en(RamSpWf_en),
    .addr(RamSpWf_addr),
    .di(RamSpWf_di),
    .dout(RamSpWf_dout)
  );
  assign io_dataRead = RamSpWf_dout; // @[Memory.scala 63:17]
  assign RamSpWf_clk = clock; // @[Memory.scala 58:21]
  assign RamSpWf_we = io_writeEnable; // @[Memory.scala 59:20]
  assign RamSpWf_en = 1'h1; // @[Memory.scala 60:20]
  assign RamSpWf_addr = io_address; // @[Memory.scala 61:22]
  assign RamSpWf_di = io_dataWrite; // @[Memory.scala 62:20]
endmodule
module Memory_34(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [10:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5), .LOAD_FILE("memory_init/backbuffer_init.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 5'h0; // @[Memory.scala 70:20]
endmodule
module Memory_35(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_36(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_37(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_38(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_39(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_40(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_41(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_42(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_43(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_8.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_44(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_9.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_45(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_10.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_46(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_11.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_47(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_12.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_48(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_13.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_49(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_14.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_50(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_15.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module MultiHotPriortyReductionTree(
  input  [5:0] io_dataInput_0,
  input  [5:0] io_dataInput_1,
  input  [5:0] io_dataInput_2,
  input  [5:0] io_dataInput_3,
  input  [5:0] io_dataInput_4,
  input  [5:0] io_dataInput_5,
  input  [5:0] io_dataInput_6,
  input  [5:0] io_dataInput_7,
  input  [5:0] io_dataInput_8,
  input  [5:0] io_dataInput_9,
  input  [5:0] io_dataInput_10,
  input  [5:0] io_dataInput_11,
  input  [5:0] io_dataInput_12,
  input  [5:0] io_dataInput_13,
  input  [5:0] io_dataInput_14,
  input  [5:0] io_dataInput_15,
  input        io_selectInput_0,
  input        io_selectInput_1,
  input        io_selectInput_2,
  input        io_selectInput_3,
  input        io_selectInput_4,
  input        io_selectInput_5,
  input        io_selectInput_6,
  input        io_selectInput_7,
  input        io_selectInput_8,
  input        io_selectInput_9,
  input        io_selectInput_10,
  input        io_selectInput_11,
  input        io_selectInput_12,
  input        io_selectInput_13,
  input        io_selectInput_14,
  input        io_selectInput_15,
  output [5:0] io_dataOutput,
  output       io_selectOutput
);
  wire  selectNodeOutputs_7 = io_selectInput_0 | io_selectInput_1; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_8 = io_selectInput_2 | io_selectInput_3; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_3 = selectNodeOutputs_7 | selectNodeOutputs_8; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_9 = io_selectInput_4 | io_selectInput_5; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_10 = io_selectInput_6 | io_selectInput_7; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_4 = selectNodeOutputs_9 | selectNodeOutputs_10; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_1 = selectNodeOutputs_3 | selectNodeOutputs_4; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_7 = io_selectInput_0 ? io_dataInput_0 : io_dataInput_1; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_8 = io_selectInput_2 ? io_dataInput_2 : io_dataInput_3; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_3 = selectNodeOutputs_7 ? dataNodeOutputs_7 : dataNodeOutputs_8; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_9 = io_selectInput_4 ? io_dataInput_4 : io_dataInput_5; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_10 = io_selectInput_6 ? io_dataInput_6 : io_dataInput_7; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_4 = selectNodeOutputs_9 ? dataNodeOutputs_9 : dataNodeOutputs_10; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_1 = selectNodeOutputs_3 ? dataNodeOutputs_3 : dataNodeOutputs_4; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_11 = io_selectInput_8 | io_selectInput_9; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_12 = io_selectInput_10 | io_selectInput_11; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_5 = selectNodeOutputs_11 | selectNodeOutputs_12; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_11 = io_selectInput_8 ? io_dataInput_8 : io_dataInput_9; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_12 = io_selectInput_10 ? io_dataInput_10 : io_dataInput_11; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_5 = selectNodeOutputs_11 ? dataNodeOutputs_11 : dataNodeOutputs_12; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_13 = io_selectInput_12 | io_selectInput_13; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_13 = io_selectInput_12 ? io_dataInput_12 : io_dataInput_13; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_14 = io_selectInput_14 ? io_dataInput_14 : io_dataInput_15; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_6 = selectNodeOutputs_13 ? dataNodeOutputs_13 : dataNodeOutputs_14; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_2 = selectNodeOutputs_5 ? dataNodeOutputs_5 : dataNodeOutputs_6; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_14 = io_selectInput_14 | io_selectInput_15; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_6 = selectNodeOutputs_13 | selectNodeOutputs_14; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_2 = selectNodeOutputs_5 | selectNodeOutputs_6; // @[GameUtilities.scala 86:54]
  assign io_dataOutput = selectNodeOutputs_1 ? dataNodeOutputs_1 : dataNodeOutputs_2; // @[GameUtilities.scala 72:17]
  assign io_selectOutput = selectNodeOutputs_1 | selectNodeOutputs_2; // @[GameUtilities.scala 73:19]
endmodule
module GraphicEngineVGA(
  input         clock,
  input         reset,
  input  [10:0] io_spriteXPosition_0,
  input  [9:0]  io_spriteYPosition_0,
  input         io_spriteFlipHorizontal_0,
  output        io_newFrame,
  input         io_frameUpdateDone,
  output        io_missingFrameError,
  output [3:0]  io_vgaRed,
  output [3:0]  io_vgaBlue,
  output [3:0]  io_vgaGreen,
  output        io_Hsync,
  output        io_Vsync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
`endif // RANDOMIZE_REG_INIT
  wire  backTileMemories_0_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_0_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_1_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_1_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_2_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_2_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_2_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_3_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_3_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_3_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_4_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_4_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_4_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_5_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_5_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_5_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_6_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_6_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_6_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_7_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_7_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_7_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_8_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_8_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_8_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_9_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_9_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_9_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_10_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_10_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_10_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_11_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_11_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_11_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_12_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_12_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_12_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_13_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_13_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_13_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_14_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_14_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_14_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_15_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_15_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_15_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_16_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_16_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_16_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_17_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_17_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_17_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_18_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_18_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_18_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_19_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_19_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_19_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_20_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_20_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_20_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_21_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_21_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_21_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_22_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_22_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_22_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_23_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_23_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_23_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_24_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_24_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_24_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_25_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_25_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_25_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_26_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_26_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_26_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_27_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_27_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_27_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_28_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_28_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_28_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_29_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_29_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_29_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_30_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_30_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_30_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backTileMemories_31_clock; // @[GraphicEngineVGA.scala 165:32]
  wire [9:0] backTileMemories_31_io_address; // @[GraphicEngineVGA.scala 165:32]
  wire [6:0] backTileMemories_31_io_dataRead; // @[GraphicEngineVGA.scala 165:32]
  wire  backBufferMemory_clock; // @[GraphicEngineVGA.scala 182:32]
  wire [10:0] backBufferMemory_io_address; // @[GraphicEngineVGA.scala 182:32]
  wire [4:0] backBufferMemory_io_dataRead; // @[GraphicEngineVGA.scala 182:32]
  wire  backBufferMemory_io_writeEnable; // @[GraphicEngineVGA.scala 182:32]
  wire [4:0] backBufferMemory_io_dataWrite; // @[GraphicEngineVGA.scala 182:32]
  wire  backBufferShadowMemory_clock; // @[GraphicEngineVGA.scala 183:38]
  wire [10:0] backBufferShadowMemory_io_address; // @[GraphicEngineVGA.scala 183:38]
  wire [4:0] backBufferShadowMemory_io_dataRead; // @[GraphicEngineVGA.scala 183:38]
  wire  backBufferShadowMemory_io_writeEnable; // @[GraphicEngineVGA.scala 183:38]
  wire [4:0] backBufferShadowMemory_io_dataWrite; // @[GraphicEngineVGA.scala 183:38]
  wire  backBufferRestoreMemory_clock; // @[GraphicEngineVGA.scala 184:39]
  wire [10:0] backBufferRestoreMemory_io_address; // @[GraphicEngineVGA.scala 184:39]
  wire [4:0] backBufferRestoreMemory_io_dataRead; // @[GraphicEngineVGA.scala 184:39]
  wire  spriteMemories_0_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_0_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_1_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_1_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_2_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_2_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_2_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_3_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_3_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_3_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_4_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_4_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_4_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_5_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_5_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_5_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_6_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_6_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_6_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_7_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_7_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_7_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_8_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_8_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_8_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_9_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_9_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_9_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_10_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_10_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_10_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_11_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_11_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_11_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_12_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_12_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_12_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_13_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_13_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_13_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_14_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_14_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_14_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire  spriteMemories_15_clock; // @[GraphicEngineVGA.scala 254:30]
  wire [9:0] spriteMemories_15_io_address; // @[GraphicEngineVGA.scala 254:30]
  wire [6:0] spriteMemories_15_io_dataRead; // @[GraphicEngineVGA.scala 254:30]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_0; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_1; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_2; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_3; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_4; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_5; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_6; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_7; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_8; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_9; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_10; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_11; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_12; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_13; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_14; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_15; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_0; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_1; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_2; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_3; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_4; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_5; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_6; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_7; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_8; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_9; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_10; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_11; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_12; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_13; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_14; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectInput_15; // @[GraphicEngineVGA.scala 372:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataOutput; // @[GraphicEngineVGA.scala 372:44]
  wire  multiHotPriortyReductionTree_io_selectOutput; // @[GraphicEngineVGA.scala 372:44]
  reg [1:0] ScaleCounterReg; // @[GraphicEngineVGA.scala 68:32]
  reg [9:0] CounterXReg; // @[GraphicEngineVGA.scala 69:28]
  reg [9:0] CounterYReg; // @[GraphicEngineVGA.scala 70:28]
  wire  _T = ScaleCounterReg == 2'h3; // @[GraphicEngineVGA.scala 76:26]
  wire  _T_1 = CounterXReg == 10'h31f; // @[GraphicEngineVGA.scala 79:24]
  wire  _T_2 = CounterYReg == 10'h20c; // @[GraphicEngineVGA.scala 81:26]
  wire [9:0] _T_4 = CounterYReg + 10'h1; // @[GraphicEngineVGA.scala 85:38]
  wire [9:0] _T_6 = CounterXReg + 10'h1; // @[GraphicEngineVGA.scala 88:36]
  wire  _GEN_4 = _T_1 & _T_2; // @[GraphicEngineVGA.scala 79:129]
  wire [1:0] _T_8 = ScaleCounterReg + 2'h1; // @[GraphicEngineVGA.scala 91:42]
  wire  _GEN_8 = _T & _GEN_4; // @[GraphicEngineVGA.scala 76:52]
  reg [11:0] backMemoryRestoreCounter; // @[GraphicEngineVGA.scala 206:41]
  wire  restoreEnabled = backMemoryRestoreCounter < 12'h800; // @[GraphicEngineVGA.scala 209:33]
  wire  run = restoreEnabled ? 1'h0 : 1'h1; // @[GraphicEngineVGA.scala 209:70]
  wire  _T_9 = CounterXReg >= 10'h290; // @[GraphicEngineVGA.scala 95:28]
  wire  _T_10 = CounterXReg < 10'h2f0; // @[GraphicEngineVGA.scala 95:95]
  wire  Hsync = _T_9 & _T_10; // @[GraphicEngineVGA.scala 95:79]
  wire  _T_11 = CounterYReg >= 10'h1ea; // @[GraphicEngineVGA.scala 96:28]
  wire  _T_12 = CounterYReg < 10'h1ec; // @[GraphicEngineVGA.scala 96:95]
  wire  Vsync = _T_11 & _T_12; // @[GraphicEngineVGA.scala 96:79]
  reg  _T_14_0; // @[GameUtilities.scala 21:24]
  reg  _T_14_1; // @[GameUtilities.scala 21:24]
  reg  _T_14_2; // @[GameUtilities.scala 21:24]
  reg  _T_14_3; // @[GameUtilities.scala 21:24]
  reg  _T_16_0; // @[GameUtilities.scala 21:24]
  reg  _T_16_1; // @[GameUtilities.scala 21:24]
  reg  _T_16_2; // @[GameUtilities.scala 21:24]
  reg  _T_16_3; // @[GameUtilities.scala 21:24]
  wire  _T_17 = CounterXReg < 10'h280; // @[GraphicEngineVGA.scala 100:36]
  wire  _T_18 = CounterYReg < 10'h1e0; // @[GraphicEngineVGA.scala 100:76]
  reg [20:0] frameClockCount; // @[GraphicEngineVGA.scala 107:32]
  wire  _T_19 = frameClockCount == 21'h19a27f; // @[GraphicEngineVGA.scala 108:42]
  wire [20:0] _T_21 = frameClockCount + 21'h1; // @[GraphicEngineVGA.scala 108:92]
  wire  preDisplayArea = frameClockCount >= 21'h199a1b; // @[GraphicEngineVGA.scala 109:40]
  reg [10:0] spriteXPositionReg_0; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_1; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_2; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_3; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_4; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_5; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_6; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_0; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_1; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_2; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_3; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_4; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_5; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_6; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_7; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_8; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_9; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_10; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_11; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_12; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_13; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_14; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_15; // @[Reg.scala 27:20]
  wire  _GEN_52 = io_newFrame ? 1'h0 : spriteVisibleReg_7; // @[Reg.scala 28:19]
  wire  _GEN_53 = io_newFrame ? 1'h0 : spriteVisibleReg_8; // @[Reg.scala 28:19]
  wire  _GEN_54 = io_newFrame ? 1'h0 : spriteVisibleReg_9; // @[Reg.scala 28:19]
  wire  _GEN_55 = io_newFrame ? 1'h0 : spriteVisibleReg_10; // @[Reg.scala 28:19]
  wire  _GEN_56 = io_newFrame ? 1'h0 : spriteVisibleReg_11; // @[Reg.scala 28:19]
  wire  _GEN_57 = io_newFrame ? 1'h0 : spriteVisibleReg_12; // @[Reg.scala 28:19]
  wire  _GEN_58 = io_newFrame ? 1'h0 : spriteVisibleReg_13; // @[Reg.scala 28:19]
  wire  _GEN_59 = io_newFrame ? 1'h0 : spriteVisibleReg_14; // @[Reg.scala 28:19]
  wire  _GEN_60 = io_newFrame ? 1'h0 : spriteVisibleReg_15; // @[Reg.scala 28:19]
  reg  spriteFlipHorizontalReg_0; // @[Reg.scala 27:20]
  reg  spriteFlipHorizontalReg_1; // @[Reg.scala 27:20]
  reg  spriteFlipHorizontalReg_4; // @[Reg.scala 27:20]
  wire  _GEN_62 = io_newFrame | spriteFlipHorizontalReg_1; // @[Reg.scala 28:19]
  wire  _GEN_65 = io_newFrame | spriteFlipHorizontalReg_4; // @[Reg.scala 28:19]
  reg  spriteFlipVerticalReg_2; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_5; // @[Reg.scala 27:20]
  wire  _GEN_79 = io_newFrame | spriteFlipVerticalReg_2; // @[Reg.scala 28:19]
  wire  _GEN_82 = io_newFrame | spriteFlipVerticalReg_5; // @[Reg.scala 28:19]
  reg [1:0] spriteScaleHorizontalReg_0; // @[Reg.scala 27:20]
  reg [1:0] spriteScaleHorizontalReg_1; // @[Reg.scala 27:20]
  reg [1:0] spriteScaleHorizontalReg_2; // @[Reg.scala 27:20]
  reg [1:0] spriteScaleHorizontalReg_4; // @[Reg.scala 27:20]
  reg [1:0] spriteScaleVerticalReg_0; // @[Reg.scala 27:20]
  reg [1:0] spriteScaleVerticalReg_1; // @[Reg.scala 27:20]
  reg [1:0] spriteScaleVerticalReg_2; // @[Reg.scala 27:20]
  reg [1:0] spriteScaleVerticalReg_4; // @[Reg.scala 27:20]
  reg  spriteRotationReg_4; // @[Reg.scala 27:20]
  reg  spriteRotationReg_6; // @[Reg.scala 27:20]
  wire  _GEN_129 = io_newFrame | spriteRotationReg_4; // @[Reg.scala 28:19]
  wire  _GEN_131 = io_newFrame | spriteRotationReg_6; // @[Reg.scala 28:19]
  reg  missingFrameErrorReg; // @[GraphicEngineVGA.scala 132:37]
  wire [10:0] pixelXBack = {{1'd0}, CounterXReg}; // @[GraphicEngineVGA.scala 143:27]
  wire [10:0] pixelYBack = {{1'd0}, CounterYReg}; // @[GraphicEngineVGA.scala 144:27]
  reg  newFrameStikyReg; // @[GraphicEngineVGA.scala 151:33]
  wire  _GEN_144 = io_newFrame | newFrameStikyReg; // @[GraphicEngineVGA.scala 152:21]
  reg  _T_36; // @[GraphicEngineVGA.scala 155:15]
  wire  _T_37 = newFrameStikyReg & io_newFrame; // @[GraphicEngineVGA.scala 158:25]
  wire  _GEN_146 = _T_37 | missingFrameErrorReg; // @[GraphicEngineVGA.scala 158:41]
  wire [5:0] _GEN_67900 = {{1'd0}, pixelYBack[4:0]}; // @[GraphicEngineVGA.scala 176:76]
  wire [10:0] _T_40 = 6'h20 * _GEN_67900; // @[GraphicEngineVGA.scala 176:76]
  wire [10:0] _GEN_67901 = {{6'd0}, pixelXBack[4:0]}; // @[GraphicEngineVGA.scala 176:63]
  wire [11:0] _T_41 = _GEN_67901 + _T_40; // @[GraphicEngineVGA.scala 176:63]
  reg [6:0] backTileMemoryDataRead_0; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_1; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_2; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_3; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_4; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_5; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_6; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_7; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_8; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_9; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_10; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_11; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_12; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_13; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_14; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_15; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_16; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_17; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_18; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_19; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_20; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_21; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_22; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_23; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_24; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_25; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_26; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_27; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_28; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_29; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_30; // @[GraphicEngineVGA.scala 177:41]
  reg [6:0] backTileMemoryDataRead_31; // @[GraphicEngineVGA.scala 177:41]
  reg [11:0] backMemoryCopyCounter; // @[GraphicEngineVGA.scala 187:38]
  wire  _T_198 = backMemoryCopyCounter < 12'h800; // @[GraphicEngineVGA.scala 191:32]
  wire [11:0] _T_200 = backMemoryCopyCounter + 12'h1; // @[GraphicEngineVGA.scala 192:54]
  wire  copyEnabled = preDisplayArea & _T_198; // @[GraphicEngineVGA.scala 190:24]
  reg  copyEnabledReg; // @[GraphicEngineVGA.scala 204:31]
  wire [11:0] _T_203 = backMemoryRestoreCounter + 12'h1; // @[GraphicEngineVGA.scala 210:58]
  reg [10:0] _T_206; // @[GraphicEngineVGA.scala 225:67]
  wire [10:0] _T_209 = copyEnabled ? backMemoryCopyCounter[10:0] : 11'h0; // @[GraphicEngineVGA.scala 225:105]
  reg  _T_211; // @[GraphicEngineVGA.scala 227:71]
  reg [10:0] _T_218; // @[GraphicEngineVGA.scala 230:61]
  wire [11:0] _T_221 = 6'h28 * pixelYBack[10:5]; // @[GraphicEngineVGA.scala 230:131]
  wire [11:0] _GEN_67964 = {{6'd0}, pixelXBack[10:5]}; // @[GraphicEngineVGA.scala 230:118]
  wire [12:0] _T_222 = _GEN_67964 + _T_221; // @[GraphicEngineVGA.scala 230:118]
  wire [12:0] _T_223 = copyEnabledReg ? {{2'd0}, _T_218} : _T_222; // @[GraphicEngineVGA.scala 230:37]
  reg [4:0] _T_225; // @[GraphicEngineVGA.scala 247:56]
  wire [6:0] _GEN_157 = 5'h1 == _T_225 ? backTileMemoryDataRead_1 : backTileMemoryDataRead_0; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_158 = 5'h2 == _T_225 ? backTileMemoryDataRead_2 : _GEN_157; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_159 = 5'h3 == _T_225 ? backTileMemoryDataRead_3 : _GEN_158; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_160 = 5'h4 == _T_225 ? backTileMemoryDataRead_4 : _GEN_159; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_161 = 5'h5 == _T_225 ? backTileMemoryDataRead_5 : _GEN_160; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_162 = 5'h6 == _T_225 ? backTileMemoryDataRead_6 : _GEN_161; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_163 = 5'h7 == _T_225 ? backTileMemoryDataRead_7 : _GEN_162; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_164 = 5'h8 == _T_225 ? backTileMemoryDataRead_8 : _GEN_163; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_165 = 5'h9 == _T_225 ? backTileMemoryDataRead_9 : _GEN_164; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_166 = 5'ha == _T_225 ? backTileMemoryDataRead_10 : _GEN_165; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_167 = 5'hb == _T_225 ? backTileMemoryDataRead_11 : _GEN_166; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_168 = 5'hc == _T_225 ? backTileMemoryDataRead_12 : _GEN_167; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_169 = 5'hd == _T_225 ? backTileMemoryDataRead_13 : _GEN_168; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_170 = 5'he == _T_225 ? backTileMemoryDataRead_14 : _GEN_169; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_171 = 5'hf == _T_225 ? backTileMemoryDataRead_15 : _GEN_170; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_172 = 5'h10 == _T_225 ? backTileMemoryDataRead_16 : _GEN_171; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_173 = 5'h11 == _T_225 ? backTileMemoryDataRead_17 : _GEN_172; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_174 = 5'h12 == _T_225 ? backTileMemoryDataRead_18 : _GEN_173; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_175 = 5'h13 == _T_225 ? backTileMemoryDataRead_19 : _GEN_174; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_176 = 5'h14 == _T_225 ? backTileMemoryDataRead_20 : _GEN_175; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_177 = 5'h15 == _T_225 ? backTileMemoryDataRead_21 : _GEN_176; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_178 = 5'h16 == _T_225 ? backTileMemoryDataRead_22 : _GEN_177; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_179 = 5'h17 == _T_225 ? backTileMemoryDataRead_23 : _GEN_178; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_180 = 5'h18 == _T_225 ? backTileMemoryDataRead_24 : _GEN_179; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_181 = 5'h19 == _T_225 ? backTileMemoryDataRead_25 : _GEN_180; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_182 = 5'h1a == _T_225 ? backTileMemoryDataRead_26 : _GEN_181; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_183 = 5'h1b == _T_225 ? backTileMemoryDataRead_27 : _GEN_182; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_184 = 5'h1c == _T_225 ? backTileMemoryDataRead_28 : _GEN_183; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_185 = 5'h1d == _T_225 ? backTileMemoryDataRead_29 : _GEN_184; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] _GEN_186 = 5'h1e == _T_225 ? backTileMemoryDataRead_30 : _GEN_185; // @[GraphicEngineVGA.scala 247:23]
  wire [6:0] fullBackgroundColor = 5'h1f == _T_225 ? backTileMemoryDataRead_31 : _GEN_186; // @[GraphicEngineVGA.scala 247:23]
  reg [5:0] pixelColorBack; // @[GraphicEngineVGA.scala 249:31]
  wire [10:0] _T_232 = {1'h0,CounterXReg}; // @[GraphicEngineVGA.scala 301:66]
  wire [11:0] _T_233 = $signed(_T_232) - $signed(spriteXPositionReg_0); // @[GraphicEngineVGA.scala 301:73]
  wire [10:0] _T_242 = {1'h0,CounterYReg}; // @[GraphicEngineVGA.scala 302:66]
  wire [10:0] _GEN_67965 = {{1{spriteYPositionReg_0[9]}},spriteYPositionReg_0}; // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_243 = $signed(_T_242) - $signed(_GEN_67965); // @[GraphicEngineVGA.scala 302:73]
  wire  _T_258 = 2'h2 == spriteScaleHorizontalReg_0; // @[Mux.scala 80:60]
  wire [7:0] _T_259 = _T_258 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_260 = 2'h1 == spriteScaleHorizontalReg_0; // @[Mux.scala 80:60]
  wire [7:0] _T_261 = _T_260 ? $signed(8'sh10) : $signed(_T_259); // @[Mux.scala 80:57]
  wire  _T_262 = 2'h0 == spriteScaleHorizontalReg_0; // @[Mux.scala 80:60]
  wire [7:0] _T_263 = _T_262 ? $signed(8'sh20) : $signed(_T_261); // @[Mux.scala 80:57]
  wire  _T_264 = 2'h2 == spriteScaleVerticalReg_0; // @[Mux.scala 80:60]
  wire [7:0] _T_265 = _T_264 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_266 = 2'h1 == spriteScaleVerticalReg_0; // @[Mux.scala 80:60]
  wire [7:0] _T_267 = _T_266 ? $signed(8'sh10) : $signed(_T_265); // @[Mux.scala 80:57]
  wire  _T_268 = 2'h0 == spriteScaleVerticalReg_0; // @[Mux.scala 80:60]
  wire [7:0] _T_269 = _T_268 ? $signed(8'sh20) : $signed(_T_267); // @[Mux.scala 80:57]
  wire [7:0] _T_272 = $signed(_T_263) - 8'sh1; // @[GraphicEngineVGA.scala 338:58]
  wire [11:0] _GEN_67968 = {{4{_T_272[7]}},_T_272}; // @[GraphicEngineVGA.scala 338:65]
  wire [11:0] _T_275 = $signed(_GEN_67968) - $signed(_T_233); // @[GraphicEngineVGA.scala 338:65]
  wire [11:0] _T_276 = spriteFlipHorizontalReg_0 ? $signed(_T_275) : $signed(_T_233); // @[GraphicEngineVGA.scala 338:23]
  wire [10:0] inSpriteY_0 = _T_243[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire  _T_291 = $signed(_T_276) >= 12'sh0; // @[GraphicEngineVGA.scala 347:31]
  wire [11:0] _GEN_67971 = {{4{_T_263[7]}},_T_263}; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_292 = $signed(_T_276) < $signed(_GEN_67971); // @[GraphicEngineVGA.scala 347:52]
  wire  _T_293 = _T_291 & _T_292; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_294 = $signed(inSpriteY_0) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire [10:0] _GEN_67972 = {{3{_T_269[7]}},_T_269}; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_295 = $signed(inSpriteY_0) < $signed(_GEN_67972); // @[GraphicEngineVGA.scala 348:52]
  wire  _T_296 = _T_294 & _T_295; // @[GraphicEngineVGA.scala 348:39]
  wire [10:0] _T_302 = _T_276[11:1]; // @[GraphicEngineVGA.scala 354:24]
  wire [6:0] _T_305 = _T_276[4:0] * 5'h2; // @[GraphicEngineVGA.scala 355:36]
  wire [4:0] _T_308 = _T_258 ? _T_302[4:0] : _T_276[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_310 = _T_260 ? _T_305 : {{2'd0}, _T_308}; // @[Mux.scala 80:57]
  wire [6:0] _T_312 = _T_262 ? {{2'd0}, _T_276[4:0]} : _T_310; // @[Mux.scala 80:57]
  wire [9:0] _T_314 = inSpriteY_0[10:1]; // @[GraphicEngineVGA.scala 359:24]
  wire [6:0] _T_317 = inSpriteY_0[4:0] * 5'h2; // @[GraphicEngineVGA.scala 360:36]
  wire [4:0] _T_320 = _T_264 ? _T_314[4:0] : inSpriteY_0[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_322 = _T_266 ? _T_317 : {{2'd0}, _T_320}; // @[Mux.scala 80:57]
  wire [6:0] _T_324 = _T_268 ? {{2'd0}, inSpriteY_0[4:0]} : _T_322; // @[Mux.scala 80:57]
  wire [12:0] _T_325 = 7'h20 * _T_324; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_67973 = {{6'd0}, _T_312}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_327 = _GEN_67973 + _T_325; // @[GraphicEngineVGA.scala 367:46]
  wire [11:0] _T_330 = $signed(_T_232) - $signed(spriteXPositionReg_1); // @[GraphicEngineVGA.scala 301:73]
  wire [10:0] _GEN_67974 = {{1{spriteYPositionReg_1[9]}},spriteYPositionReg_1}; // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_340 = $signed(_T_242) - $signed(_GEN_67974); // @[GraphicEngineVGA.scala 302:73]
  wire  _T_355 = 2'h2 == spriteScaleHorizontalReg_1; // @[Mux.scala 80:60]
  wire [7:0] _T_356 = _T_355 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_357 = 2'h1 == spriteScaleHorizontalReg_1; // @[Mux.scala 80:60]
  wire [7:0] _T_358 = _T_357 ? $signed(8'sh10) : $signed(_T_356); // @[Mux.scala 80:57]
  wire  _T_359 = 2'h0 == spriteScaleHorizontalReg_1; // @[Mux.scala 80:60]
  wire [7:0] _T_360 = _T_359 ? $signed(8'sh20) : $signed(_T_358); // @[Mux.scala 80:57]
  wire  _T_361 = 2'h2 == spriteScaleVerticalReg_1; // @[Mux.scala 80:60]
  wire [7:0] _T_362 = _T_361 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_363 = 2'h1 == spriteScaleVerticalReg_1; // @[Mux.scala 80:60]
  wire [7:0] _T_364 = _T_363 ? $signed(8'sh10) : $signed(_T_362); // @[Mux.scala 80:57]
  wire  _T_365 = 2'h0 == spriteScaleVerticalReg_1; // @[Mux.scala 80:60]
  wire [7:0] _T_366 = _T_365 ? $signed(8'sh20) : $signed(_T_364); // @[Mux.scala 80:57]
  wire [7:0] _T_369 = $signed(_T_360) - 8'sh1; // @[GraphicEngineVGA.scala 338:58]
  wire [11:0] _GEN_67977 = {{4{_T_369[7]}},_T_369}; // @[GraphicEngineVGA.scala 338:65]
  wire [11:0] _T_372 = $signed(_GEN_67977) - $signed(_T_330); // @[GraphicEngineVGA.scala 338:65]
  wire [11:0] _T_373 = spriteFlipHorizontalReg_1 ? $signed(_T_372) : $signed(_T_330); // @[GraphicEngineVGA.scala 338:23]
  wire [10:0] inSpriteY_1 = _T_340[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire  _T_388 = $signed(_T_373) >= 12'sh0; // @[GraphicEngineVGA.scala 347:31]
  wire [11:0] _GEN_67980 = {{4{_T_360[7]}},_T_360}; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_389 = $signed(_T_373) < $signed(_GEN_67980); // @[GraphicEngineVGA.scala 347:52]
  wire  _T_390 = _T_388 & _T_389; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_391 = $signed(inSpriteY_1) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire [10:0] _GEN_67981 = {{3{_T_366[7]}},_T_366}; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_392 = $signed(inSpriteY_1) < $signed(_GEN_67981); // @[GraphicEngineVGA.scala 348:52]
  wire  _T_393 = _T_391 & _T_392; // @[GraphicEngineVGA.scala 348:39]
  wire [10:0] _T_399 = _T_373[11:1]; // @[GraphicEngineVGA.scala 354:24]
  wire [6:0] _T_402 = _T_373[4:0] * 5'h2; // @[GraphicEngineVGA.scala 355:36]
  wire [4:0] _T_405 = _T_355 ? _T_399[4:0] : _T_373[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_407 = _T_357 ? _T_402 : {{2'd0}, _T_405}; // @[Mux.scala 80:57]
  wire [6:0] _T_409 = _T_359 ? {{2'd0}, _T_373[4:0]} : _T_407; // @[Mux.scala 80:57]
  wire [9:0] _T_411 = inSpriteY_1[10:1]; // @[GraphicEngineVGA.scala 359:24]
  wire [6:0] _T_414 = inSpriteY_1[4:0] * 5'h2; // @[GraphicEngineVGA.scala 360:36]
  wire [4:0] _T_417 = _T_361 ? _T_411[4:0] : inSpriteY_1[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_419 = _T_363 ? _T_414 : {{2'd0}, _T_417}; // @[Mux.scala 80:57]
  wire [6:0] _T_421 = _T_365 ? {{2'd0}, inSpriteY_1[4:0]} : _T_419; // @[Mux.scala 80:57]
  wire [12:0] _T_422 = 7'h20 * _T_421; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_67982 = {{6'd0}, _T_409}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_424 = _GEN_67982 + _T_422; // @[GraphicEngineVGA.scala 367:46]
  wire [11:0] _T_427 = $signed(_T_232) - $signed(spriteXPositionReg_2); // @[GraphicEngineVGA.scala 301:73]
  wire [10:0] _GEN_67983 = {{1{spriteYPositionReg_2[9]}},spriteYPositionReg_2}; // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_437 = $signed(_T_242) - $signed(_GEN_67983); // @[GraphicEngineVGA.scala 302:73]
  wire  _T_452 = 2'h2 == spriteScaleHorizontalReg_2; // @[Mux.scala 80:60]
  wire [7:0] _T_453 = _T_452 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_454 = 2'h1 == spriteScaleHorizontalReg_2; // @[Mux.scala 80:60]
  wire [7:0] _T_455 = _T_454 ? $signed(8'sh10) : $signed(_T_453); // @[Mux.scala 80:57]
  wire  _T_456 = 2'h0 == spriteScaleHorizontalReg_2; // @[Mux.scala 80:60]
  wire [7:0] _T_457 = _T_456 ? $signed(8'sh20) : $signed(_T_455); // @[Mux.scala 80:57]
  wire  _T_458 = 2'h2 == spriteScaleVerticalReg_2; // @[Mux.scala 80:60]
  wire [7:0] _T_459 = _T_458 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_460 = 2'h1 == spriteScaleVerticalReg_2; // @[Mux.scala 80:60]
  wire [7:0] _T_461 = _T_460 ? $signed(8'sh10) : $signed(_T_459); // @[Mux.scala 80:57]
  wire  _T_462 = 2'h0 == spriteScaleVerticalReg_2; // @[Mux.scala 80:60]
  wire [7:0] _T_463 = _T_462 ? $signed(8'sh20) : $signed(_T_461); // @[Mux.scala 80:57]
  wire [7:0] _T_473 = $signed(_T_463) - 8'sh1; // @[GraphicEngineVGA.scala 339:58]
  wire [10:0] inSpriteY_2 = _T_437[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire [10:0] _GEN_67988 = {{3{_T_473[7]}},_T_473}; // @[GraphicEngineVGA.scala 339:65]
  wire [10:0] _T_476 = $signed(_GEN_67988) - $signed(inSpriteY_2); // @[GraphicEngineVGA.scala 339:65]
  wire [10:0] _T_477 = spriteFlipVerticalReg_2 ? $signed(_T_476) : $signed(inSpriteY_2); // @[GraphicEngineVGA.scala 339:23]
  wire  _T_478 = $signed(_T_427) >= 12'sh0; // @[GraphicEngineVGA.scala 343:27]
  wire [11:0] _GEN_67989 = {{4{_T_457[7]}},_T_457}; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_486 = $signed(_T_427) < $signed(_GEN_67989); // @[GraphicEngineVGA.scala 347:52]
  wire  _T_487 = _T_478 & _T_486; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_488 = $signed(_T_477) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire [10:0] _GEN_67990 = {{3{_T_463[7]}},_T_463}; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_489 = $signed(_T_477) < $signed(_GEN_67990); // @[GraphicEngineVGA.scala 348:52]
  wire  _T_490 = _T_488 & _T_489; // @[GraphicEngineVGA.scala 348:39]
  wire [10:0] _T_496 = _T_427[11:1]; // @[GraphicEngineVGA.scala 354:24]
  wire [6:0] _T_499 = _T_427[4:0] * 5'h2; // @[GraphicEngineVGA.scala 355:36]
  wire [4:0] _T_502 = _T_452 ? _T_496[4:0] : _T_427[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_504 = _T_454 ? _T_499 : {{2'd0}, _T_502}; // @[Mux.scala 80:57]
  wire [6:0] _T_506 = _T_456 ? {{2'd0}, _T_427[4:0]} : _T_504; // @[Mux.scala 80:57]
  wire [9:0] _T_508 = _T_477[10:1]; // @[GraphicEngineVGA.scala 359:24]
  wire [6:0] _T_511 = _T_477[4:0] * 5'h2; // @[GraphicEngineVGA.scala 360:36]
  wire [4:0] _T_514 = _T_458 ? _T_508[4:0] : _T_477[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_516 = _T_460 ? _T_511 : {{2'd0}, _T_514}; // @[Mux.scala 80:57]
  wire [6:0] _T_518 = _T_462 ? {{2'd0}, _T_477[4:0]} : _T_516; // @[Mux.scala 80:57]
  wire [12:0] _T_519 = 7'h20 * _T_518; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_67991 = {{6'd0}, _T_506}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_521 = _GEN_67991 + _T_519; // @[GraphicEngineVGA.scala 367:46]
  wire [11:0] _T_524 = $signed(_T_232) - $signed(spriteXPositionReg_3); // @[GraphicEngineVGA.scala 301:73]
  wire [10:0] _GEN_67992 = {{1{spriteYPositionReg_3[9]}},spriteYPositionReg_3}; // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_534 = $signed(_T_242) - $signed(_GEN_67992); // @[GraphicEngineVGA.scala 302:73]
  wire [7:0] _T_563 = 8'sh20 - 8'sh1; // @[GraphicEngineVGA.scala 338:58]
  wire [10:0] inSpriteY_3 = _T_534[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire [10:0] _GEN_67997 = {{3{_T_563[7]}},_T_563}; // @[GraphicEngineVGA.scala 339:65]
  wire  _T_575 = $signed(_T_524) >= 12'sh0; // @[GraphicEngineVGA.scala 343:27]
  wire  _T_583 = $signed(_T_524) < 12'sh20; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_584 = _T_575 & _T_583; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_585 = $signed(inSpriteY_3) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire  _T_586 = $signed(inSpriteY_3) < 11'sh20; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_587 = _T_585 & _T_586; // @[GraphicEngineVGA.scala 348:39]
  wire [6:0] _T_601 = {{2'd0}, _T_524[4:0]}; // @[Mux.scala 80:57]
  wire [6:0] _T_613 = {{2'd0}, inSpriteY_3[4:0]}; // @[Mux.scala 80:57]
  wire [12:0] _T_616 = 7'h20 * _T_613; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_67998 = {{6'd0}, _T_601}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_618 = _GEN_67998 + _T_616; // @[GraphicEngineVGA.scala 367:46]
  wire [11:0] _T_621 = $signed(_T_232) - $signed(spriteXPositionReg_4); // @[GraphicEngineVGA.scala 301:73]
  wire [11:0] _T_624 = $signed(_T_621) + 12'sh7; // @[GraphicEngineVGA.scala 301:98]
  wire [11:0] _T_628 = spriteRotationReg_4 ? $signed(_T_624) : $signed(_T_621); // @[GraphicEngineVGA.scala 301:22]
  wire [10:0] _GEN_67999 = {{1{spriteYPositionReg_4[9]}},spriteYPositionReg_4}; // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_631 = $signed(_T_242) - $signed(_GEN_67999); // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_634 = $signed(_T_631) + 12'sh7; // @[GraphicEngineVGA.scala 302:98]
  wire [11:0] _T_638 = spriteRotationReg_4 ? $signed(_T_634) : $signed(_T_631); // @[GraphicEngineVGA.scala 302:22]
  wire [11:0] _T_640 = _T_638[5:0] * 6'h2e; // @[GraphicEngineVGA.scala 307:34]
  wire [11:0] _GEN_68001 = {{6'd0}, _T_628[5:0]}; // @[GraphicEngineVGA.scala 307:53]
  wire [11:0] _T_643 = _T_640 + _GEN_68001; // @[GraphicEngineVGA.scala 307:53]
  wire [6:0] _GEN_17117 = 12'h1 == _T_643 ? $signed(-7'sh10) : $signed(-7'sh11); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17118 = 12'h2 == _T_643 ? $signed(-7'shf) : $signed(_GEN_17117); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17119 = 12'h3 == _T_643 ? $signed(-7'she) : $signed(_GEN_17118); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17120 = 12'h4 == _T_643 ? $signed(-7'she) : $signed(_GEN_17119); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17121 = 12'h5 == _T_643 ? $signed(-7'shd) : $signed(_GEN_17120); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17122 = 12'h6 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17121); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17123 = 12'h7 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17122); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17124 = 12'h8 == _T_643 ? $signed(-7'shb) : $signed(_GEN_17123); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17125 = 12'h9 == _T_643 ? $signed(-7'sha) : $signed(_GEN_17124); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17126 = 12'ha == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17125); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17127 = 12'hb == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17126); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17128 = 12'hc == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17127); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17129 = 12'hd == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17128); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17130 = 12'he == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17129); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17131 = 12'hf == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17130); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17132 = 12'h10 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17131); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17133 = 12'h11 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17132); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17134 = 12'h12 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17133); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17135 = 12'h13 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17134); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17136 = 12'h14 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17135); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17137 = 12'h15 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17136); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17138 = 12'h16 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17137); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17139 = 12'h17 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17138); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17140 = 12'h18 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17139); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17141 = 12'h19 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17140); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17142 = 12'h1a == _T_643 ? $signed(7'sh2) : $signed(_GEN_17141); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17143 = 12'h1b == _T_643 ? $signed(7'sh3) : $signed(_GEN_17142); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17144 = 12'h1c == _T_643 ? $signed(7'sh3) : $signed(_GEN_17143); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17145 = 12'h1d == _T_643 ? $signed(7'sh4) : $signed(_GEN_17144); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17146 = 12'h1e == _T_643 ? $signed(7'sh5) : $signed(_GEN_17145); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17147 = 12'h1f == _T_643 ? $signed(7'sh5) : $signed(_GEN_17146); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17148 = 12'h20 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17147); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17149 = 12'h21 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17148); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17150 = 12'h22 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17149); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17151 = 12'h23 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17150); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17152 = 12'h24 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17151); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17153 = 12'h25 == _T_643 ? $signed(7'sha) : $signed(_GEN_17152); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17154 = 12'h26 == _T_643 ? $signed(7'sha) : $signed(_GEN_17153); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17155 = 12'h27 == _T_643 ? $signed(7'shb) : $signed(_GEN_17154); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17156 = 12'h28 == _T_643 ? $signed(7'shc) : $signed(_GEN_17155); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17157 = 12'h29 == _T_643 ? $signed(7'shc) : $signed(_GEN_17156); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17158 = 12'h2a == _T_643 ? $signed(7'shd) : $signed(_GEN_17157); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17159 = 12'h2b == _T_643 ? $signed(7'she) : $signed(_GEN_17158); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17160 = 12'h2c == _T_643 ? $signed(7'shf) : $signed(_GEN_17159); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17161 = 12'h2d == _T_643 ? $signed(7'shf) : $signed(_GEN_17160); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17162 = 12'h2e == _T_643 ? $signed(-7'sh10) : $signed(_GEN_17161); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17163 = 12'h2f == _T_643 ? $signed(-7'shf) : $signed(_GEN_17162); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17164 = 12'h30 == _T_643 ? $signed(-7'she) : $signed(_GEN_17163); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17165 = 12'h31 == _T_643 ? $signed(-7'she) : $signed(_GEN_17164); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17166 = 12'h32 == _T_643 ? $signed(-7'shd) : $signed(_GEN_17165); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17167 = 12'h33 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17166); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17168 = 12'h34 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17167); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17169 = 12'h35 == _T_643 ? $signed(-7'shb) : $signed(_GEN_17168); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17170 = 12'h36 == _T_643 ? $signed(-7'sha) : $signed(_GEN_17169); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17171 = 12'h37 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17170); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17172 = 12'h38 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17171); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17173 = 12'h39 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17172); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17174 = 12'h3a == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17173); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17175 = 12'h3b == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17174); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17176 = 12'h3c == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17175); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17177 = 12'h3d == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17176); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17178 = 12'h3e == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17177); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17179 = 12'h3f == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17178); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17180 = 12'h40 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17179); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17181 = 12'h41 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17180); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17182 = 12'h42 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17181); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17183 = 12'h43 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17182); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17184 = 12'h44 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17183); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17185 = 12'h45 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17184); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17186 = 12'h46 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17185); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17187 = 12'h47 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17186); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17188 = 12'h48 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17187); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17189 = 12'h49 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17188); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17190 = 12'h4a == _T_643 ? $signed(7'sh4) : $signed(_GEN_17189); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17191 = 12'h4b == _T_643 ? $signed(7'sh5) : $signed(_GEN_17190); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17192 = 12'h4c == _T_643 ? $signed(7'sh5) : $signed(_GEN_17191); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17193 = 12'h4d == _T_643 ? $signed(7'sh6) : $signed(_GEN_17192); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17194 = 12'h4e == _T_643 ? $signed(7'sh7) : $signed(_GEN_17193); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17195 = 12'h4f == _T_643 ? $signed(7'sh8) : $signed(_GEN_17194); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17196 = 12'h50 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17195); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17197 = 12'h51 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17196); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17198 = 12'h52 == _T_643 ? $signed(7'sha) : $signed(_GEN_17197); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17199 = 12'h53 == _T_643 ? $signed(7'sha) : $signed(_GEN_17198); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17200 = 12'h54 == _T_643 ? $signed(7'shb) : $signed(_GEN_17199); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17201 = 12'h55 == _T_643 ? $signed(7'shc) : $signed(_GEN_17200); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17202 = 12'h56 == _T_643 ? $signed(7'shc) : $signed(_GEN_17201); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17203 = 12'h57 == _T_643 ? $signed(7'shd) : $signed(_GEN_17202); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17204 = 12'h58 == _T_643 ? $signed(7'she) : $signed(_GEN_17203); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17205 = 12'h59 == _T_643 ? $signed(7'shf) : $signed(_GEN_17204); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17206 = 12'h5a == _T_643 ? $signed(7'shf) : $signed(_GEN_17205); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17207 = 12'h5b == _T_643 ? $signed(7'sh10) : $signed(_GEN_17206); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17208 = 12'h5c == _T_643 ? $signed(-7'shf) : $signed(_GEN_17207); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17209 = 12'h5d == _T_643 ? $signed(-7'she) : $signed(_GEN_17208); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17210 = 12'h5e == _T_643 ? $signed(-7'she) : $signed(_GEN_17209); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17211 = 12'h5f == _T_643 ? $signed(-7'shd) : $signed(_GEN_17210); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17212 = 12'h60 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17211); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17213 = 12'h61 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17212); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17214 = 12'h62 == _T_643 ? $signed(-7'shb) : $signed(_GEN_17213); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17215 = 12'h63 == _T_643 ? $signed(-7'sha) : $signed(_GEN_17214); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17216 = 12'h64 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17215); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17217 = 12'h65 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17216); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17218 = 12'h66 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17217); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17219 = 12'h67 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17218); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17220 = 12'h68 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17219); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17221 = 12'h69 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17220); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17222 = 12'h6a == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17221); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17223 = 12'h6b == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17222); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17224 = 12'h6c == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17223); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17225 = 12'h6d == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17224); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17226 = 12'h6e == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17225); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17227 = 12'h6f == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17226); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17228 = 12'h70 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17227); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17229 = 12'h71 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17228); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17230 = 12'h72 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17229); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17231 = 12'h73 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17230); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17232 = 12'h74 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17231); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17233 = 12'h75 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17232); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17234 = 12'h76 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17233); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17235 = 12'h77 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17234); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17236 = 12'h78 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17235); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17237 = 12'h79 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17236); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17238 = 12'h7a == _T_643 ? $signed(7'sh6) : $signed(_GEN_17237); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17239 = 12'h7b == _T_643 ? $signed(7'sh7) : $signed(_GEN_17238); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17240 = 12'h7c == _T_643 ? $signed(7'sh8) : $signed(_GEN_17239); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17241 = 12'h7d == _T_643 ? $signed(7'sh8) : $signed(_GEN_17240); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17242 = 12'h7e == _T_643 ? $signed(7'sh9) : $signed(_GEN_17241); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17243 = 12'h7f == _T_643 ? $signed(7'sha) : $signed(_GEN_17242); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17244 = 12'h80 == _T_643 ? $signed(7'sha) : $signed(_GEN_17243); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17245 = 12'h81 == _T_643 ? $signed(7'shb) : $signed(_GEN_17244); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17246 = 12'h82 == _T_643 ? $signed(7'shc) : $signed(_GEN_17245); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17247 = 12'h83 == _T_643 ? $signed(7'shc) : $signed(_GEN_17246); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17248 = 12'h84 == _T_643 ? $signed(7'shd) : $signed(_GEN_17247); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17249 = 12'h85 == _T_643 ? $signed(7'she) : $signed(_GEN_17248); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17250 = 12'h86 == _T_643 ? $signed(7'shf) : $signed(_GEN_17249); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17251 = 12'h87 == _T_643 ? $signed(7'shf) : $signed(_GEN_17250); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17252 = 12'h88 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17251); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17253 = 12'h89 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17252); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17254 = 12'h8a == _T_643 ? $signed(-7'she) : $signed(_GEN_17253); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17255 = 12'h8b == _T_643 ? $signed(-7'she) : $signed(_GEN_17254); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17256 = 12'h8c == _T_643 ? $signed(-7'shd) : $signed(_GEN_17255); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17257 = 12'h8d == _T_643 ? $signed(-7'shc) : $signed(_GEN_17256); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17258 = 12'h8e == _T_643 ? $signed(-7'shc) : $signed(_GEN_17257); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17259 = 12'h8f == _T_643 ? $signed(-7'shb) : $signed(_GEN_17258); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17260 = 12'h90 == _T_643 ? $signed(-7'sha) : $signed(_GEN_17259); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17261 = 12'h91 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17260); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17262 = 12'h92 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17261); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17263 = 12'h93 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17262); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17264 = 12'h94 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17263); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17265 = 12'h95 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17264); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17266 = 12'h96 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17265); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17267 = 12'h97 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17266); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17268 = 12'h98 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17267); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17269 = 12'h99 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17268); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17270 = 12'h9a == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17269); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17271 = 12'h9b == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17270); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17272 = 12'h9c == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17271); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17273 = 12'h9d == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17272); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17274 = 12'h9e == _T_643 ? $signed(7'sh0) : $signed(_GEN_17273); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17275 = 12'h9f == _T_643 ? $signed(7'sh0) : $signed(_GEN_17274); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17276 = 12'ha0 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17275); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17277 = 12'ha1 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17276); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17278 = 12'ha2 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17277); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17279 = 12'ha3 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17278); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17280 = 12'ha4 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17279); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17281 = 12'ha5 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17280); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17282 = 12'ha6 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17281); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17283 = 12'ha7 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17282); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17284 = 12'ha8 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17283); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17285 = 12'ha9 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17284); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17286 = 12'haa == _T_643 ? $signed(7'sh8) : $signed(_GEN_17285); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17287 = 12'hab == _T_643 ? $signed(7'sh9) : $signed(_GEN_17286); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17288 = 12'hac == _T_643 ? $signed(7'sha) : $signed(_GEN_17287); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17289 = 12'had == _T_643 ? $signed(7'sha) : $signed(_GEN_17288); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17290 = 12'hae == _T_643 ? $signed(7'shb) : $signed(_GEN_17289); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17291 = 12'haf == _T_643 ? $signed(7'shc) : $signed(_GEN_17290); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17292 = 12'hb0 == _T_643 ? $signed(7'shc) : $signed(_GEN_17291); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17293 = 12'hb1 == _T_643 ? $signed(7'shd) : $signed(_GEN_17292); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17294 = 12'hb2 == _T_643 ? $signed(7'she) : $signed(_GEN_17293); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17295 = 12'hb3 == _T_643 ? $signed(7'shf) : $signed(_GEN_17294); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17296 = 12'hb4 == _T_643 ? $signed(7'shf) : $signed(_GEN_17295); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17297 = 12'hb5 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17296); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17298 = 12'hb6 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17297); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17299 = 12'hb7 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17298); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17300 = 12'hb8 == _T_643 ? $signed(-7'she) : $signed(_GEN_17299); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17301 = 12'hb9 == _T_643 ? $signed(-7'shd) : $signed(_GEN_17300); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17302 = 12'hba == _T_643 ? $signed(-7'shc) : $signed(_GEN_17301); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17303 = 12'hbb == _T_643 ? $signed(-7'shc) : $signed(_GEN_17302); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17304 = 12'hbc == _T_643 ? $signed(-7'shb) : $signed(_GEN_17303); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17305 = 12'hbd == _T_643 ? $signed(-7'sha) : $signed(_GEN_17304); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17306 = 12'hbe == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17305); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17307 = 12'hbf == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17306); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17308 = 12'hc0 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17307); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17309 = 12'hc1 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17308); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17310 = 12'hc2 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17309); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17311 = 12'hc3 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17310); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17312 = 12'hc4 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17311); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17313 = 12'hc5 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17312); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17314 = 12'hc6 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17313); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17315 = 12'hc7 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17314); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17316 = 12'hc8 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17315); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17317 = 12'hc9 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17316); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17318 = 12'hca == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17317); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17319 = 12'hcb == _T_643 ? $signed(7'sh0) : $signed(_GEN_17318); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17320 = 12'hcc == _T_643 ? $signed(7'sh0) : $signed(_GEN_17319); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17321 = 12'hcd == _T_643 ? $signed(7'sh1) : $signed(_GEN_17320); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17322 = 12'hce == _T_643 ? $signed(7'sh2) : $signed(_GEN_17321); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17323 = 12'hcf == _T_643 ? $signed(7'sh3) : $signed(_GEN_17322); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17324 = 12'hd0 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17323); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17325 = 12'hd1 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17324); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17326 = 12'hd2 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17325); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17327 = 12'hd3 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17326); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17328 = 12'hd4 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17327); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17329 = 12'hd5 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17328); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17330 = 12'hd6 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17329); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17331 = 12'hd7 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17330); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17332 = 12'hd8 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17331); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17333 = 12'hd9 == _T_643 ? $signed(7'sha) : $signed(_GEN_17332); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17334 = 12'hda == _T_643 ? $signed(7'sha) : $signed(_GEN_17333); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17335 = 12'hdb == _T_643 ? $signed(7'shb) : $signed(_GEN_17334); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17336 = 12'hdc == _T_643 ? $signed(7'shc) : $signed(_GEN_17335); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17337 = 12'hdd == _T_643 ? $signed(7'shc) : $signed(_GEN_17336); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17338 = 12'hde == _T_643 ? $signed(7'shd) : $signed(_GEN_17337); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17339 = 12'hdf == _T_643 ? $signed(7'she) : $signed(_GEN_17338); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17340 = 12'he0 == _T_643 ? $signed(7'shf) : $signed(_GEN_17339); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17341 = 12'he1 == _T_643 ? $signed(7'shf) : $signed(_GEN_17340); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17342 = 12'he2 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17341); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17343 = 12'he3 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17342); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17344 = 12'he4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17343); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17345 = 12'he5 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17344); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17346 = 12'he6 == _T_643 ? $signed(-7'shd) : $signed(_GEN_17345); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17347 = 12'he7 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17346); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17348 = 12'he8 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17347); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17349 = 12'he9 == _T_643 ? $signed(-7'shb) : $signed(_GEN_17348); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17350 = 12'hea == _T_643 ? $signed(-7'sha) : $signed(_GEN_17349); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17351 = 12'heb == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17350); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17352 = 12'hec == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17351); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17353 = 12'hed == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17352); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17354 = 12'hee == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17353); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17355 = 12'hef == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17354); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17356 = 12'hf0 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17355); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17357 = 12'hf1 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17356); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17358 = 12'hf2 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17357); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17359 = 12'hf3 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17358); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17360 = 12'hf4 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17359); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17361 = 12'hf5 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17360); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17362 = 12'hf6 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17361); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17363 = 12'hf7 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17362); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17364 = 12'hf8 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17363); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17365 = 12'hf9 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17364); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17366 = 12'hfa == _T_643 ? $signed(7'sh1) : $signed(_GEN_17365); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17367 = 12'hfb == _T_643 ? $signed(7'sh2) : $signed(_GEN_17366); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17368 = 12'hfc == _T_643 ? $signed(7'sh3) : $signed(_GEN_17367); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17369 = 12'hfd == _T_643 ? $signed(7'sh3) : $signed(_GEN_17368); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17370 = 12'hfe == _T_643 ? $signed(7'sh4) : $signed(_GEN_17369); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17371 = 12'hff == _T_643 ? $signed(7'sh5) : $signed(_GEN_17370); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17372 = 12'h100 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17371); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17373 = 12'h101 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17372); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17374 = 12'h102 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17373); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17375 = 12'h103 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17374); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17376 = 12'h104 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17375); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17377 = 12'h105 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17376); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17378 = 12'h106 == _T_643 ? $signed(7'sha) : $signed(_GEN_17377); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17379 = 12'h107 == _T_643 ? $signed(7'sha) : $signed(_GEN_17378); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17380 = 12'h108 == _T_643 ? $signed(7'shb) : $signed(_GEN_17379); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17381 = 12'h109 == _T_643 ? $signed(7'shc) : $signed(_GEN_17380); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17382 = 12'h10a == _T_643 ? $signed(7'shc) : $signed(_GEN_17381); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17383 = 12'h10b == _T_643 ? $signed(7'shd) : $signed(_GEN_17382); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17384 = 12'h10c == _T_643 ? $signed(7'she) : $signed(_GEN_17383); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17385 = 12'h10d == _T_643 ? $signed(7'shf) : $signed(_GEN_17384); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17386 = 12'h10e == _T_643 ? $signed(7'shf) : $signed(_GEN_17385); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17387 = 12'h10f == _T_643 ? $signed(7'sh10) : $signed(_GEN_17386); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17388 = 12'h110 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17387); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17389 = 12'h111 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17388); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17390 = 12'h112 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17389); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17391 = 12'h113 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17390); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17392 = 12'h114 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17391); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17393 = 12'h115 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17392); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17394 = 12'h116 == _T_643 ? $signed(-7'shb) : $signed(_GEN_17393); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17395 = 12'h117 == _T_643 ? $signed(-7'sha) : $signed(_GEN_17394); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17396 = 12'h118 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17395); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17397 = 12'h119 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17396); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17398 = 12'h11a == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17397); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17399 = 12'h11b == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17398); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17400 = 12'h11c == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17399); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17401 = 12'h11d == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17400); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17402 = 12'h11e == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17401); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17403 = 12'h11f == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17402); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17404 = 12'h120 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17403); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17405 = 12'h121 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17404); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17406 = 12'h122 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17405); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17407 = 12'h123 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17406); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17408 = 12'h124 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17407); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17409 = 12'h125 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17408); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17410 = 12'h126 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17409); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17411 = 12'h127 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17410); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17412 = 12'h128 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17411); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17413 = 12'h129 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17412); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17414 = 12'h12a == _T_643 ? $signed(7'sh3) : $signed(_GEN_17413); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17415 = 12'h12b == _T_643 ? $signed(7'sh4) : $signed(_GEN_17414); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17416 = 12'h12c == _T_643 ? $signed(7'sh5) : $signed(_GEN_17415); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17417 = 12'h12d == _T_643 ? $signed(7'sh5) : $signed(_GEN_17416); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17418 = 12'h12e == _T_643 ? $signed(7'sh6) : $signed(_GEN_17417); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17419 = 12'h12f == _T_643 ? $signed(7'sh7) : $signed(_GEN_17418); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17420 = 12'h130 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17419); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17421 = 12'h131 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17420); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17422 = 12'h132 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17421); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17423 = 12'h133 == _T_643 ? $signed(7'sha) : $signed(_GEN_17422); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17424 = 12'h134 == _T_643 ? $signed(7'sha) : $signed(_GEN_17423); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17425 = 12'h135 == _T_643 ? $signed(7'shb) : $signed(_GEN_17424); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17426 = 12'h136 == _T_643 ? $signed(7'shc) : $signed(_GEN_17425); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17427 = 12'h137 == _T_643 ? $signed(7'shc) : $signed(_GEN_17426); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17428 = 12'h138 == _T_643 ? $signed(7'shd) : $signed(_GEN_17427); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17429 = 12'h139 == _T_643 ? $signed(7'she) : $signed(_GEN_17428); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17430 = 12'h13a == _T_643 ? $signed(7'shf) : $signed(_GEN_17429); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17431 = 12'h13b == _T_643 ? $signed(7'shf) : $signed(_GEN_17430); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17432 = 12'h13c == _T_643 ? $signed(7'sh10) : $signed(_GEN_17431); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17433 = 12'h13d == _T_643 ? $signed(7'sh11) : $signed(_GEN_17432); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17434 = 12'h13e == _T_643 ? $signed(7'sh11) : $signed(_GEN_17433); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17435 = 12'h13f == _T_643 ? $signed(7'sh12) : $signed(_GEN_17434); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17436 = 12'h140 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17435); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17437 = 12'h141 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17436); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17438 = 12'h142 == _T_643 ? $signed(-7'shc) : $signed(_GEN_17437); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17439 = 12'h143 == _T_643 ? $signed(-7'shb) : $signed(_GEN_17438); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17440 = 12'h144 == _T_643 ? $signed(-7'sha) : $signed(_GEN_17439); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17441 = 12'h145 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17440); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17442 = 12'h146 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17441); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17443 = 12'h147 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17442); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17444 = 12'h148 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17443); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17445 = 12'h149 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17444); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17446 = 12'h14a == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17445); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17447 = 12'h14b == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17446); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17448 = 12'h14c == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17447); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17449 = 12'h14d == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17448); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17450 = 12'h14e == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17449); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17451 = 12'h14f == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17450); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17452 = 12'h150 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17451); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17453 = 12'h151 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17452); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17454 = 12'h152 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17453); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17455 = 12'h153 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17454); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17456 = 12'h154 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17455); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17457 = 12'h155 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17456); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17458 = 12'h156 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17457); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17459 = 12'h157 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17458); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17460 = 12'h158 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17459); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17461 = 12'h159 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17460); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17462 = 12'h15a == _T_643 ? $signed(7'sh5) : $signed(_GEN_17461); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17463 = 12'h15b == _T_643 ? $signed(7'sh6) : $signed(_GEN_17462); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17464 = 12'h15c == _T_643 ? $signed(7'sh7) : $signed(_GEN_17463); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17465 = 12'h15d == _T_643 ? $signed(7'sh8) : $signed(_GEN_17464); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17466 = 12'h15e == _T_643 ? $signed(7'sh8) : $signed(_GEN_17465); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17467 = 12'h15f == _T_643 ? $signed(7'sh9) : $signed(_GEN_17466); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17468 = 12'h160 == _T_643 ? $signed(7'sha) : $signed(_GEN_17467); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17469 = 12'h161 == _T_643 ? $signed(7'sha) : $signed(_GEN_17468); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17470 = 12'h162 == _T_643 ? $signed(7'shb) : $signed(_GEN_17469); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17471 = 12'h163 == _T_643 ? $signed(7'shc) : $signed(_GEN_17470); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17472 = 12'h164 == _T_643 ? $signed(7'shc) : $signed(_GEN_17471); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17473 = 12'h165 == _T_643 ? $signed(7'shd) : $signed(_GEN_17472); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17474 = 12'h166 == _T_643 ? $signed(7'she) : $signed(_GEN_17473); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17475 = 12'h167 == _T_643 ? $signed(7'shf) : $signed(_GEN_17474); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17476 = 12'h168 == _T_643 ? $signed(7'shf) : $signed(_GEN_17475); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17477 = 12'h169 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17476); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17478 = 12'h16a == _T_643 ? $signed(7'sh11) : $signed(_GEN_17477); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17479 = 12'h16b == _T_643 ? $signed(7'sh11) : $signed(_GEN_17478); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17480 = 12'h16c == _T_643 ? $signed(7'sh12) : $signed(_GEN_17479); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17481 = 12'h16d == _T_643 ? $signed(7'sh13) : $signed(_GEN_17480); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17482 = 12'h16e == _T_643 ? $signed(7'sh14) : $signed(_GEN_17481); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17483 = 12'h16f == _T_643 ? $signed(7'sh14) : $signed(_GEN_17482); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17484 = 12'h170 == _T_643 ? $signed(-7'shb) : $signed(_GEN_17483); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17485 = 12'h171 == _T_643 ? $signed(-7'sha) : $signed(_GEN_17484); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17486 = 12'h172 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17485); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17487 = 12'h173 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17486); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17488 = 12'h174 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17487); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17489 = 12'h175 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17488); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17490 = 12'h176 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17489); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17491 = 12'h177 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17490); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17492 = 12'h178 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17491); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17493 = 12'h179 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17492); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17494 = 12'h17a == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17493); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17495 = 12'h17b == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17494); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17496 = 12'h17c == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17495); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17497 = 12'h17d == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17496); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17498 = 12'h17e == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17497); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17499 = 12'h17f == _T_643 ? $signed(7'sh0) : $signed(_GEN_17498); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17500 = 12'h180 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17499); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17501 = 12'h181 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17500); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17502 = 12'h182 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17501); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17503 = 12'h183 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17502); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17504 = 12'h184 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17503); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17505 = 12'h185 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17504); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17506 = 12'h186 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17505); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17507 = 12'h187 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17506); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17508 = 12'h188 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17507); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17509 = 12'h189 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17508); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17510 = 12'h18a == _T_643 ? $signed(7'sh8) : $signed(_GEN_17509); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17511 = 12'h18b == _T_643 ? $signed(7'sh8) : $signed(_GEN_17510); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17512 = 12'h18c == _T_643 ? $signed(7'sh9) : $signed(_GEN_17511); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17513 = 12'h18d == _T_643 ? $signed(7'sha) : $signed(_GEN_17512); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17514 = 12'h18e == _T_643 ? $signed(7'sha) : $signed(_GEN_17513); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17515 = 12'h18f == _T_643 ? $signed(7'shb) : $signed(_GEN_17514); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17516 = 12'h190 == _T_643 ? $signed(7'shc) : $signed(_GEN_17515); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17517 = 12'h191 == _T_643 ? $signed(7'shc) : $signed(_GEN_17516); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17518 = 12'h192 == _T_643 ? $signed(7'shd) : $signed(_GEN_17517); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17519 = 12'h193 == _T_643 ? $signed(7'she) : $signed(_GEN_17518); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17520 = 12'h194 == _T_643 ? $signed(7'shf) : $signed(_GEN_17519); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17521 = 12'h195 == _T_643 ? $signed(7'shf) : $signed(_GEN_17520); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17522 = 12'h196 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17521); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17523 = 12'h197 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17522); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17524 = 12'h198 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17523); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17525 = 12'h199 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17524); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17526 = 12'h19a == _T_643 ? $signed(7'sh13) : $signed(_GEN_17525); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17527 = 12'h19b == _T_643 ? $signed(7'sh14) : $signed(_GEN_17526); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17528 = 12'h19c == _T_643 ? $signed(7'sh14) : $signed(_GEN_17527); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17529 = 12'h19d == _T_643 ? $signed(7'sh15) : $signed(_GEN_17528); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17530 = 12'h19e == _T_643 ? $signed(-7'sha) : $signed(_GEN_17529); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17531 = 12'h19f == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17530); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17532 = 12'h1a0 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17531); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17533 = 12'h1a1 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17532); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17534 = 12'h1a2 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17533); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17535 = 12'h1a3 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17534); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17536 = 12'h1a4 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17535); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17537 = 12'h1a5 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17536); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17538 = 12'h1a6 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17537); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17539 = 12'h1a7 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17538); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17540 = 12'h1a8 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17539); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17541 = 12'h1a9 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17540); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17542 = 12'h1aa == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17541); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17543 = 12'h1ab == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17542); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17544 = 12'h1ac == _T_643 ? $signed(7'sh0) : $signed(_GEN_17543); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17545 = 12'h1ad == _T_643 ? $signed(7'sh0) : $signed(_GEN_17544); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17546 = 12'h1ae == _T_643 ? $signed(7'sh1) : $signed(_GEN_17545); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17547 = 12'h1af == _T_643 ? $signed(7'sh2) : $signed(_GEN_17546); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17548 = 12'h1b0 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17547); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17549 = 12'h1b1 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17548); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17550 = 12'h1b2 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17549); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17551 = 12'h1b3 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17550); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17552 = 12'h1b4 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17551); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17553 = 12'h1b5 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17552); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17554 = 12'h1b6 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17553); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17555 = 12'h1b7 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17554); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17556 = 12'h1b8 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17555); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17557 = 12'h1b9 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17556); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17558 = 12'h1ba == _T_643 ? $signed(7'sha) : $signed(_GEN_17557); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17559 = 12'h1bb == _T_643 ? $signed(7'sha) : $signed(_GEN_17558); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17560 = 12'h1bc == _T_643 ? $signed(7'shb) : $signed(_GEN_17559); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17561 = 12'h1bd == _T_643 ? $signed(7'shc) : $signed(_GEN_17560); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17562 = 12'h1be == _T_643 ? $signed(7'shc) : $signed(_GEN_17561); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17563 = 12'h1bf == _T_643 ? $signed(7'shd) : $signed(_GEN_17562); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17564 = 12'h1c0 == _T_643 ? $signed(7'she) : $signed(_GEN_17563); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17565 = 12'h1c1 == _T_643 ? $signed(7'shf) : $signed(_GEN_17564); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17566 = 12'h1c2 == _T_643 ? $signed(7'shf) : $signed(_GEN_17565); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17567 = 12'h1c3 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17566); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17568 = 12'h1c4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17567); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17569 = 12'h1c5 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17568); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17570 = 12'h1c6 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17569); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17571 = 12'h1c7 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17570); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17572 = 12'h1c8 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17571); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17573 = 12'h1c9 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17572); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17574 = 12'h1ca == _T_643 ? $signed(7'sh15) : $signed(_GEN_17573); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17575 = 12'h1cb == _T_643 ? $signed(7'sh16) : $signed(_GEN_17574); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17576 = 12'h1cc == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17575); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17577 = 12'h1cd == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17576); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17578 = 12'h1ce == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17577); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17579 = 12'h1cf == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17578); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17580 = 12'h1d0 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17579); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17581 = 12'h1d1 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17580); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17582 = 12'h1d2 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17581); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17583 = 12'h1d3 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17582); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17584 = 12'h1d4 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17583); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17585 = 12'h1d5 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17584); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17586 = 12'h1d6 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17585); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17587 = 12'h1d7 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17586); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17588 = 12'h1d8 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17587); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17589 = 12'h1d9 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17588); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17590 = 12'h1da == _T_643 ? $signed(7'sh0) : $signed(_GEN_17589); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17591 = 12'h1db == _T_643 ? $signed(7'sh1) : $signed(_GEN_17590); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17592 = 12'h1dc == _T_643 ? $signed(7'sh2) : $signed(_GEN_17591); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17593 = 12'h1dd == _T_643 ? $signed(7'sh3) : $signed(_GEN_17592); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17594 = 12'h1de == _T_643 ? $signed(7'sh3) : $signed(_GEN_17593); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17595 = 12'h1df == _T_643 ? $signed(7'sh4) : $signed(_GEN_17594); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17596 = 12'h1e0 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17595); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17597 = 12'h1e1 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17596); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17598 = 12'h1e2 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17597); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17599 = 12'h1e3 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17598); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17600 = 12'h1e4 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17599); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17601 = 12'h1e5 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17600); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17602 = 12'h1e6 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17601); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17603 = 12'h1e7 == _T_643 ? $signed(7'sha) : $signed(_GEN_17602); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17604 = 12'h1e8 == _T_643 ? $signed(7'sha) : $signed(_GEN_17603); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17605 = 12'h1e9 == _T_643 ? $signed(7'shb) : $signed(_GEN_17604); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17606 = 12'h1ea == _T_643 ? $signed(7'shc) : $signed(_GEN_17605); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17607 = 12'h1eb == _T_643 ? $signed(7'shc) : $signed(_GEN_17606); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17608 = 12'h1ec == _T_643 ? $signed(7'shd) : $signed(_GEN_17607); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17609 = 12'h1ed == _T_643 ? $signed(7'she) : $signed(_GEN_17608); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17610 = 12'h1ee == _T_643 ? $signed(7'shf) : $signed(_GEN_17609); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17611 = 12'h1ef == _T_643 ? $signed(7'shf) : $signed(_GEN_17610); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17612 = 12'h1f0 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17611); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17613 = 12'h1f1 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17612); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17614 = 12'h1f2 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17613); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17615 = 12'h1f3 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17614); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17616 = 12'h1f4 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17615); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17617 = 12'h1f5 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17616); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17618 = 12'h1f6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17617); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17619 = 12'h1f7 == _T_643 ? $signed(7'sh15) : $signed(_GEN_17618); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17620 = 12'h1f8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17619); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17621 = 12'h1f9 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17620); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17622 = 12'h1fa == _T_643 ? $signed(-7'sh9) : $signed(_GEN_17621); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17623 = 12'h1fb == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17622); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17624 = 12'h1fc == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17623); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17625 = 12'h1fd == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17624); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17626 = 12'h1fe == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17625); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17627 = 12'h1ff == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17626); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17628 = 12'h200 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17627); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17629 = 12'h201 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17628); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17630 = 12'h202 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17629); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17631 = 12'h203 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17630); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17632 = 12'h204 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17631); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17633 = 12'h205 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17632); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17634 = 12'h206 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17633); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17635 = 12'h207 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17634); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17636 = 12'h208 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17635); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17637 = 12'h209 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17636); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17638 = 12'h20a == _T_643 ? $signed(7'sh3) : $signed(_GEN_17637); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17639 = 12'h20b == _T_643 ? $signed(7'sh3) : $signed(_GEN_17638); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17640 = 12'h20c == _T_643 ? $signed(7'sh4) : $signed(_GEN_17639); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17641 = 12'h20d == _T_643 ? $signed(7'sh5) : $signed(_GEN_17640); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17642 = 12'h20e == _T_643 ? $signed(7'sh5) : $signed(_GEN_17641); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17643 = 12'h20f == _T_643 ? $signed(7'sh6) : $signed(_GEN_17642); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17644 = 12'h210 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17643); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17645 = 12'h211 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17644); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17646 = 12'h212 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17645); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17647 = 12'h213 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17646); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17648 = 12'h214 == _T_643 ? $signed(7'sha) : $signed(_GEN_17647); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17649 = 12'h215 == _T_643 ? $signed(7'sha) : $signed(_GEN_17648); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17650 = 12'h216 == _T_643 ? $signed(7'shb) : $signed(_GEN_17649); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17651 = 12'h217 == _T_643 ? $signed(7'shc) : $signed(_GEN_17650); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17652 = 12'h218 == _T_643 ? $signed(7'shc) : $signed(_GEN_17651); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17653 = 12'h219 == _T_643 ? $signed(7'shd) : $signed(_GEN_17652); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17654 = 12'h21a == _T_643 ? $signed(7'she) : $signed(_GEN_17653); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17655 = 12'h21b == _T_643 ? $signed(7'shf) : $signed(_GEN_17654); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17656 = 12'h21c == _T_643 ? $signed(7'shf) : $signed(_GEN_17655); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17657 = 12'h21d == _T_643 ? $signed(7'sh10) : $signed(_GEN_17656); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17658 = 12'h21e == _T_643 ? $signed(7'sh11) : $signed(_GEN_17657); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17659 = 12'h21f == _T_643 ? $signed(7'sh11) : $signed(_GEN_17658); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17660 = 12'h220 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17659); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17661 = 12'h221 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17660); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17662 = 12'h222 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17661); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17663 = 12'h223 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17662); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17664 = 12'h224 == _T_643 ? $signed(7'sh15) : $signed(_GEN_17663); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17665 = 12'h225 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17664); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17666 = 12'h226 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17665); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17667 = 12'h227 == _T_643 ? $signed(7'sh17) : $signed(_GEN_17666); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17668 = 12'h228 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_17667); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17669 = 12'h229 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17668); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17670 = 12'h22a == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17669); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17671 = 12'h22b == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17670); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17672 = 12'h22c == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17671); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17673 = 12'h22d == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17672); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17674 = 12'h22e == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17673); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17675 = 12'h22f == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17674); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17676 = 12'h230 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17675); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17677 = 12'h231 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17676); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17678 = 12'h232 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17677); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17679 = 12'h233 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17678); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17680 = 12'h234 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17679); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17681 = 12'h235 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17680); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17682 = 12'h236 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17681); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17683 = 12'h237 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17682); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17684 = 12'h238 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17683); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17685 = 12'h239 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17684); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17686 = 12'h23a == _T_643 ? $signed(7'sh5) : $signed(_GEN_17685); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17687 = 12'h23b == _T_643 ? $signed(7'sh5) : $signed(_GEN_17686); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17688 = 12'h23c == _T_643 ? $signed(7'sh6) : $signed(_GEN_17687); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17689 = 12'h23d == _T_643 ? $signed(7'sh7) : $signed(_GEN_17688); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17690 = 12'h23e == _T_643 ? $signed(7'sh8) : $signed(_GEN_17689); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17691 = 12'h23f == _T_643 ? $signed(7'sh8) : $signed(_GEN_17690); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17692 = 12'h240 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17691); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17693 = 12'h241 == _T_643 ? $signed(7'sha) : $signed(_GEN_17692); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17694 = 12'h242 == _T_643 ? $signed(7'sha) : $signed(_GEN_17693); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17695 = 12'h243 == _T_643 ? $signed(7'shb) : $signed(_GEN_17694); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17696 = 12'h244 == _T_643 ? $signed(7'shc) : $signed(_GEN_17695); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17697 = 12'h245 == _T_643 ? $signed(7'shc) : $signed(_GEN_17696); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17698 = 12'h246 == _T_643 ? $signed(7'shd) : $signed(_GEN_17697); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17699 = 12'h247 == _T_643 ? $signed(7'she) : $signed(_GEN_17698); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17700 = 12'h248 == _T_643 ? $signed(7'shf) : $signed(_GEN_17699); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17701 = 12'h249 == _T_643 ? $signed(7'shf) : $signed(_GEN_17700); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17702 = 12'h24a == _T_643 ? $signed(7'sh10) : $signed(_GEN_17701); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17703 = 12'h24b == _T_643 ? $signed(7'sh11) : $signed(_GEN_17702); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17704 = 12'h24c == _T_643 ? $signed(7'sh11) : $signed(_GEN_17703); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17705 = 12'h24d == _T_643 ? $signed(7'sh12) : $signed(_GEN_17704); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17706 = 12'h24e == _T_643 ? $signed(7'sh13) : $signed(_GEN_17705); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17707 = 12'h24f == _T_643 ? $signed(7'sh14) : $signed(_GEN_17706); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17708 = 12'h250 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17707); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17709 = 12'h251 == _T_643 ? $signed(7'sh15) : $signed(_GEN_17708); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17710 = 12'h252 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17709); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17711 = 12'h253 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17710); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17712 = 12'h254 == _T_643 ? $signed(7'sh17) : $signed(_GEN_17711); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17713 = 12'h255 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17712); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17714 = 12'h256 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17713); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17715 = 12'h257 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17714); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17716 = 12'h258 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17715); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17717 = 12'h259 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17716); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17718 = 12'h25a == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17717); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17719 = 12'h25b == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17718); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17720 = 12'h25c == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17719); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17721 = 12'h25d == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17720); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17722 = 12'h25e == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17721); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17723 = 12'h25f == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17722); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17724 = 12'h260 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17723); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17725 = 12'h261 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17724); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17726 = 12'h262 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17725); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17727 = 12'h263 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17726); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17728 = 12'h264 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17727); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17729 = 12'h265 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17728); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17730 = 12'h266 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17729); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17731 = 12'h267 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17730); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17732 = 12'h268 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17731); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17733 = 12'h269 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17732); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17734 = 12'h26a == _T_643 ? $signed(7'sh7) : $signed(_GEN_17733); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17735 = 12'h26b == _T_643 ? $signed(7'sh8) : $signed(_GEN_17734); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17736 = 12'h26c == _T_643 ? $signed(7'sh8) : $signed(_GEN_17735); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17737 = 12'h26d == _T_643 ? $signed(7'sh9) : $signed(_GEN_17736); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17738 = 12'h26e == _T_643 ? $signed(7'sha) : $signed(_GEN_17737); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17739 = 12'h26f == _T_643 ? $signed(7'sha) : $signed(_GEN_17738); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17740 = 12'h270 == _T_643 ? $signed(7'shb) : $signed(_GEN_17739); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17741 = 12'h271 == _T_643 ? $signed(7'shc) : $signed(_GEN_17740); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17742 = 12'h272 == _T_643 ? $signed(7'shc) : $signed(_GEN_17741); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17743 = 12'h273 == _T_643 ? $signed(7'shd) : $signed(_GEN_17742); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17744 = 12'h274 == _T_643 ? $signed(7'she) : $signed(_GEN_17743); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17745 = 12'h275 == _T_643 ? $signed(7'shf) : $signed(_GEN_17744); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17746 = 12'h276 == _T_643 ? $signed(7'shf) : $signed(_GEN_17745); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17747 = 12'h277 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17746); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17748 = 12'h278 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17747); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17749 = 12'h279 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17748); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17750 = 12'h27a == _T_643 ? $signed(7'sh12) : $signed(_GEN_17749); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17751 = 12'h27b == _T_643 ? $signed(7'sh13) : $signed(_GEN_17750); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17752 = 12'h27c == _T_643 ? $signed(7'sh14) : $signed(_GEN_17751); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17753 = 12'h27d == _T_643 ? $signed(7'sh14) : $signed(_GEN_17752); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17754 = 12'h27e == _T_643 ? $signed(7'sh15) : $signed(_GEN_17753); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17755 = 12'h27f == _T_643 ? $signed(7'sh16) : $signed(_GEN_17754); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17756 = 12'h280 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17755); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17757 = 12'h281 == _T_643 ? $signed(7'sh17) : $signed(_GEN_17756); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17758 = 12'h282 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17757); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17759 = 12'h283 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17758); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17760 = 12'h284 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_17759); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17761 = 12'h285 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17760); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17762 = 12'h286 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17761); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17763 = 12'h287 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17762); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17764 = 12'h288 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17763); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17765 = 12'h289 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17764); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17766 = 12'h28a == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17765); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17767 = 12'h28b == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17766); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17768 = 12'h28c == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17767); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17769 = 12'h28d == _T_643 ? $signed(7'sh0) : $signed(_GEN_17768); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17770 = 12'h28e == _T_643 ? $signed(7'sh0) : $signed(_GEN_17769); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17771 = 12'h28f == _T_643 ? $signed(7'sh1) : $signed(_GEN_17770); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17772 = 12'h290 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17771); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17773 = 12'h291 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17772); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17774 = 12'h292 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17773); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17775 = 12'h293 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17774); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17776 = 12'h294 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17775); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17777 = 12'h295 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17776); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17778 = 12'h296 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17777); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17779 = 12'h297 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17778); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17780 = 12'h298 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17779); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17781 = 12'h299 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17780); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17782 = 12'h29a == _T_643 ? $signed(7'sh9) : $signed(_GEN_17781); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17783 = 12'h29b == _T_643 ? $signed(7'sha) : $signed(_GEN_17782); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17784 = 12'h29c == _T_643 ? $signed(7'sha) : $signed(_GEN_17783); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17785 = 12'h29d == _T_643 ? $signed(7'shb) : $signed(_GEN_17784); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17786 = 12'h29e == _T_643 ? $signed(7'shc) : $signed(_GEN_17785); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17787 = 12'h29f == _T_643 ? $signed(7'shc) : $signed(_GEN_17786); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17788 = 12'h2a0 == _T_643 ? $signed(7'shd) : $signed(_GEN_17787); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17789 = 12'h2a1 == _T_643 ? $signed(7'she) : $signed(_GEN_17788); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17790 = 12'h2a2 == _T_643 ? $signed(7'shf) : $signed(_GEN_17789); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17791 = 12'h2a3 == _T_643 ? $signed(7'shf) : $signed(_GEN_17790); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17792 = 12'h2a4 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17791); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17793 = 12'h2a5 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17792); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17794 = 12'h2a6 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17793); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17795 = 12'h2a7 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17794); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17796 = 12'h2a8 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17795); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17797 = 12'h2a9 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17796); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17798 = 12'h2aa == _T_643 ? $signed(7'sh14) : $signed(_GEN_17797); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17799 = 12'h2ab == _T_643 ? $signed(7'sh15) : $signed(_GEN_17798); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17800 = 12'h2ac == _T_643 ? $signed(7'sh16) : $signed(_GEN_17799); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17801 = 12'h2ad == _T_643 ? $signed(7'sh16) : $signed(_GEN_17800); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17802 = 12'h2ae == _T_643 ? $signed(7'sh17) : $signed(_GEN_17801); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17803 = 12'h2af == _T_643 ? $signed(7'sh18) : $signed(_GEN_17802); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17804 = 12'h2b0 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17803); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17805 = 12'h2b1 == _T_643 ? $signed(7'sh19) : $signed(_GEN_17804); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17806 = 12'h2b2 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_17805); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17807 = 12'h2b3 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17806); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17808 = 12'h2b4 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17807); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17809 = 12'h2b5 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17808); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17810 = 12'h2b6 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17809); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17811 = 12'h2b7 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17810); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17812 = 12'h2b8 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17811); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17813 = 12'h2b9 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17812); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17814 = 12'h2ba == _T_643 ? $signed(7'sh0) : $signed(_GEN_17813); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17815 = 12'h2bb == _T_643 ? $signed(7'sh0) : $signed(_GEN_17814); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17816 = 12'h2bc == _T_643 ? $signed(7'sh1) : $signed(_GEN_17815); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17817 = 12'h2bd == _T_643 ? $signed(7'sh2) : $signed(_GEN_17816); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17818 = 12'h2be == _T_643 ? $signed(7'sh3) : $signed(_GEN_17817); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17819 = 12'h2bf == _T_643 ? $signed(7'sh3) : $signed(_GEN_17818); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17820 = 12'h2c0 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17819); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17821 = 12'h2c1 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17820); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17822 = 12'h2c2 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17821); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17823 = 12'h2c3 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17822); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17824 = 12'h2c4 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17823); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17825 = 12'h2c5 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17824); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17826 = 12'h2c6 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17825); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17827 = 12'h2c7 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17826); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17828 = 12'h2c8 == _T_643 ? $signed(7'sha) : $signed(_GEN_17827); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17829 = 12'h2c9 == _T_643 ? $signed(7'sha) : $signed(_GEN_17828); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17830 = 12'h2ca == _T_643 ? $signed(7'shb) : $signed(_GEN_17829); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17831 = 12'h2cb == _T_643 ? $signed(7'shc) : $signed(_GEN_17830); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17832 = 12'h2cc == _T_643 ? $signed(7'shc) : $signed(_GEN_17831); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17833 = 12'h2cd == _T_643 ? $signed(7'shd) : $signed(_GEN_17832); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17834 = 12'h2ce == _T_643 ? $signed(7'she) : $signed(_GEN_17833); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17835 = 12'h2cf == _T_643 ? $signed(7'shf) : $signed(_GEN_17834); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17836 = 12'h2d0 == _T_643 ? $signed(7'shf) : $signed(_GEN_17835); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17837 = 12'h2d1 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17836); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17838 = 12'h2d2 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17837); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17839 = 12'h2d3 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17838); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17840 = 12'h2d4 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17839); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17841 = 12'h2d5 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17840); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17842 = 12'h2d6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17841); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17843 = 12'h2d7 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17842); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17844 = 12'h2d8 == _T_643 ? $signed(7'sh15) : $signed(_GEN_17843); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17845 = 12'h2d9 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17844); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17846 = 12'h2da == _T_643 ? $signed(7'sh16) : $signed(_GEN_17845); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17847 = 12'h2db == _T_643 ? $signed(7'sh17) : $signed(_GEN_17846); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17848 = 12'h2dc == _T_643 ? $signed(7'sh18) : $signed(_GEN_17847); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17849 = 12'h2dd == _T_643 ? $signed(7'sh18) : $signed(_GEN_17848); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17850 = 12'h2de == _T_643 ? $signed(7'sh19) : $signed(_GEN_17849); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17851 = 12'h2df == _T_643 ? $signed(7'sh1a) : $signed(_GEN_17850); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17852 = 12'h2e0 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17851); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17853 = 12'h2e1 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17852); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17854 = 12'h2e2 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17853); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17855 = 12'h2e3 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17854); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17856 = 12'h2e4 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17855); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17857 = 12'h2e5 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17856); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17858 = 12'h2e6 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17857); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17859 = 12'h2e7 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17858); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17860 = 12'h2e8 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17859); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17861 = 12'h2e9 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17860); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17862 = 12'h2ea == _T_643 ? $signed(7'sh2) : $signed(_GEN_17861); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17863 = 12'h2eb == _T_643 ? $signed(7'sh3) : $signed(_GEN_17862); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17864 = 12'h2ec == _T_643 ? $signed(7'sh3) : $signed(_GEN_17863); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17865 = 12'h2ed == _T_643 ? $signed(7'sh4) : $signed(_GEN_17864); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17866 = 12'h2ee == _T_643 ? $signed(7'sh5) : $signed(_GEN_17865); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17867 = 12'h2ef == _T_643 ? $signed(7'sh5) : $signed(_GEN_17866); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17868 = 12'h2f0 == _T_643 ? $signed(7'sh6) : $signed(_GEN_17867); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17869 = 12'h2f1 == _T_643 ? $signed(7'sh7) : $signed(_GEN_17868); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17870 = 12'h2f2 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17869); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17871 = 12'h2f3 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17870); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17872 = 12'h2f4 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17871); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17873 = 12'h2f5 == _T_643 ? $signed(7'sha) : $signed(_GEN_17872); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17874 = 12'h2f6 == _T_643 ? $signed(7'sha) : $signed(_GEN_17873); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17875 = 12'h2f7 == _T_643 ? $signed(7'shb) : $signed(_GEN_17874); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17876 = 12'h2f8 == _T_643 ? $signed(7'shc) : $signed(_GEN_17875); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17877 = 12'h2f9 == _T_643 ? $signed(7'shc) : $signed(_GEN_17876); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17878 = 12'h2fa == _T_643 ? $signed(7'shd) : $signed(_GEN_17877); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17879 = 12'h2fb == _T_643 ? $signed(7'she) : $signed(_GEN_17878); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17880 = 12'h2fc == _T_643 ? $signed(7'shf) : $signed(_GEN_17879); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17881 = 12'h2fd == _T_643 ? $signed(7'shf) : $signed(_GEN_17880); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17882 = 12'h2fe == _T_643 ? $signed(7'sh10) : $signed(_GEN_17881); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17883 = 12'h2ff == _T_643 ? $signed(7'sh11) : $signed(_GEN_17882); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17884 = 12'h300 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17883); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17885 = 12'h301 == _T_643 ? $signed(7'sh12) : $signed(_GEN_17884); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17886 = 12'h302 == _T_643 ? $signed(7'sh13) : $signed(_GEN_17885); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17887 = 12'h303 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17886); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17888 = 12'h304 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17887); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17889 = 12'h305 == _T_643 ? $signed(7'sh15) : $signed(_GEN_17888); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17890 = 12'h306 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17889); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17891 = 12'h307 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17890); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17892 = 12'h308 == _T_643 ? $signed(7'sh17) : $signed(_GEN_17891); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17893 = 12'h309 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17892); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17894 = 12'h30a == _T_643 ? $signed(7'sh18) : $signed(_GEN_17893); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17895 = 12'h30b == _T_643 ? $signed(7'sh19) : $signed(_GEN_17894); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17896 = 12'h30c == _T_643 ? $signed(7'sh1a) : $signed(_GEN_17895); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17897 = 12'h30d == _T_643 ? $signed(7'sh1b) : $signed(_GEN_17896); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17898 = 12'h30e == _T_643 ? $signed(-7'sh5) : $signed(_GEN_17897); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17899 = 12'h30f == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17898); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17900 = 12'h310 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17899); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17901 = 12'h311 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17900); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17902 = 12'h312 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17901); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17903 = 12'h313 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17902); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17904 = 12'h314 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17903); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17905 = 12'h315 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17904); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17906 = 12'h316 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17905); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17907 = 12'h317 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17906); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17908 = 12'h318 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17907); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17909 = 12'h319 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17908); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17910 = 12'h31a == _T_643 ? $signed(7'sh4) : $signed(_GEN_17909); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17911 = 12'h31b == _T_643 ? $signed(7'sh5) : $signed(_GEN_17910); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17912 = 12'h31c == _T_643 ? $signed(7'sh5) : $signed(_GEN_17911); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17913 = 12'h31d == _T_643 ? $signed(7'sh6) : $signed(_GEN_17912); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17914 = 12'h31e == _T_643 ? $signed(7'sh7) : $signed(_GEN_17913); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17915 = 12'h31f == _T_643 ? $signed(7'sh8) : $signed(_GEN_17914); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17916 = 12'h320 == _T_643 ? $signed(7'sh8) : $signed(_GEN_17915); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17917 = 12'h321 == _T_643 ? $signed(7'sh9) : $signed(_GEN_17916); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17918 = 12'h322 == _T_643 ? $signed(7'sha) : $signed(_GEN_17917); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17919 = 12'h323 == _T_643 ? $signed(7'sha) : $signed(_GEN_17918); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17920 = 12'h324 == _T_643 ? $signed(7'shb) : $signed(_GEN_17919); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17921 = 12'h325 == _T_643 ? $signed(7'shc) : $signed(_GEN_17920); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17922 = 12'h326 == _T_643 ? $signed(7'shc) : $signed(_GEN_17921); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17923 = 12'h327 == _T_643 ? $signed(7'shd) : $signed(_GEN_17922); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17924 = 12'h328 == _T_643 ? $signed(7'she) : $signed(_GEN_17923); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17925 = 12'h329 == _T_643 ? $signed(7'shf) : $signed(_GEN_17924); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17926 = 12'h32a == _T_643 ? $signed(7'shf) : $signed(_GEN_17925); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17927 = 12'h32b == _T_643 ? $signed(7'sh10) : $signed(_GEN_17926); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17928 = 12'h32c == _T_643 ? $signed(7'sh11) : $signed(_GEN_17927); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17929 = 12'h32d == _T_643 ? $signed(7'sh11) : $signed(_GEN_17928); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17930 = 12'h32e == _T_643 ? $signed(7'sh12) : $signed(_GEN_17929); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17931 = 12'h32f == _T_643 ? $signed(7'sh13) : $signed(_GEN_17930); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17932 = 12'h330 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17931); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17933 = 12'h331 == _T_643 ? $signed(7'sh14) : $signed(_GEN_17932); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17934 = 12'h332 == _T_643 ? $signed(7'sh15) : $signed(_GEN_17933); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17935 = 12'h333 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17934); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17936 = 12'h334 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17935); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17937 = 12'h335 == _T_643 ? $signed(7'sh17) : $signed(_GEN_17936); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17938 = 12'h336 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17937); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17939 = 12'h337 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17938); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17940 = 12'h338 == _T_643 ? $signed(7'sh19) : $signed(_GEN_17939); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17941 = 12'h339 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_17940); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17942 = 12'h33a == _T_643 ? $signed(7'sh1b) : $signed(_GEN_17941); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17943 = 12'h33b == _T_643 ? $signed(7'sh1b) : $signed(_GEN_17942); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17944 = 12'h33c == _T_643 ? $signed(-7'sh4) : $signed(_GEN_17943); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17945 = 12'h33d == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17944); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17946 = 12'h33e == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17945); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17947 = 12'h33f == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17946); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17948 = 12'h340 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17947); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17949 = 12'h341 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17948); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17950 = 12'h342 == _T_643 ? $signed(7'sh0) : $signed(_GEN_17949); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17951 = 12'h343 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17950); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17952 = 12'h344 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17951); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17953 = 12'h345 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17952); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17954 = 12'h346 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17953); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17955 = 12'h347 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17954); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17956 = 12'h348 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17955); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17957 = 12'h349 == _T_643 ? $signed(7'sh5) : $signed(_GEN_17956); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17958 = 12'h34a == _T_643 ? $signed(7'sh6) : $signed(_GEN_17957); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17959 = 12'h34b == _T_643 ? $signed(7'sh7) : $signed(_GEN_17958); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17960 = 12'h34c == _T_643 ? $signed(7'sh8) : $signed(_GEN_17959); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17961 = 12'h34d == _T_643 ? $signed(7'sh8) : $signed(_GEN_17960); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17962 = 12'h34e == _T_643 ? $signed(7'sh9) : $signed(_GEN_17961); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17963 = 12'h34f == _T_643 ? $signed(7'sha) : $signed(_GEN_17962); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17964 = 12'h350 == _T_643 ? $signed(7'sha) : $signed(_GEN_17963); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17965 = 12'h351 == _T_643 ? $signed(7'shb) : $signed(_GEN_17964); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17966 = 12'h352 == _T_643 ? $signed(7'shc) : $signed(_GEN_17965); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17967 = 12'h353 == _T_643 ? $signed(7'shc) : $signed(_GEN_17966); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17968 = 12'h354 == _T_643 ? $signed(7'shd) : $signed(_GEN_17967); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17969 = 12'h355 == _T_643 ? $signed(7'she) : $signed(_GEN_17968); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17970 = 12'h356 == _T_643 ? $signed(7'shf) : $signed(_GEN_17969); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17971 = 12'h357 == _T_643 ? $signed(7'shf) : $signed(_GEN_17970); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17972 = 12'h358 == _T_643 ? $signed(7'sh10) : $signed(_GEN_17971); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17973 = 12'h359 == _T_643 ? $signed(7'sh11) : $signed(_GEN_17972); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17974 = 12'h35a == _T_643 ? $signed(7'sh11) : $signed(_GEN_17973); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17975 = 12'h35b == _T_643 ? $signed(7'sh12) : $signed(_GEN_17974); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17976 = 12'h35c == _T_643 ? $signed(7'sh13) : $signed(_GEN_17975); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17977 = 12'h35d == _T_643 ? $signed(7'sh14) : $signed(_GEN_17976); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17978 = 12'h35e == _T_643 ? $signed(7'sh14) : $signed(_GEN_17977); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17979 = 12'h35f == _T_643 ? $signed(7'sh15) : $signed(_GEN_17978); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17980 = 12'h360 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17979); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17981 = 12'h361 == _T_643 ? $signed(7'sh16) : $signed(_GEN_17980); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17982 = 12'h362 == _T_643 ? $signed(7'sh17) : $signed(_GEN_17981); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17983 = 12'h363 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17982); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17984 = 12'h364 == _T_643 ? $signed(7'sh18) : $signed(_GEN_17983); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17985 = 12'h365 == _T_643 ? $signed(7'sh19) : $signed(_GEN_17984); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17986 = 12'h366 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_17985); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17987 = 12'h367 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_17986); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17988 = 12'h368 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_17987); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17989 = 12'h369 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_17988); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17990 = 12'h36a == _T_643 ? $signed(-7'sh3) : $signed(_GEN_17989); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17991 = 12'h36b == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17990); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17992 = 12'h36c == _T_643 ? $signed(-7'sh2) : $signed(_GEN_17991); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17993 = 12'h36d == _T_643 ? $signed(-7'sh1) : $signed(_GEN_17992); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17994 = 12'h36e == _T_643 ? $signed(7'sh0) : $signed(_GEN_17993); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17995 = 12'h36f == _T_643 ? $signed(7'sh0) : $signed(_GEN_17994); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17996 = 12'h370 == _T_643 ? $signed(7'sh1) : $signed(_GEN_17995); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17997 = 12'h371 == _T_643 ? $signed(7'sh2) : $signed(_GEN_17996); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17998 = 12'h372 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17997); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_17999 = 12'h373 == _T_643 ? $signed(7'sh3) : $signed(_GEN_17998); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18000 = 12'h374 == _T_643 ? $signed(7'sh4) : $signed(_GEN_17999); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18001 = 12'h375 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18000); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18002 = 12'h376 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18001); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18003 = 12'h377 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18002); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18004 = 12'h378 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18003); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18005 = 12'h379 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18004); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18006 = 12'h37a == _T_643 ? $signed(7'sh8) : $signed(_GEN_18005); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18007 = 12'h37b == _T_643 ? $signed(7'sh9) : $signed(_GEN_18006); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18008 = 12'h37c == _T_643 ? $signed(7'sha) : $signed(_GEN_18007); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18009 = 12'h37d == _T_643 ? $signed(7'sha) : $signed(_GEN_18008); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18010 = 12'h37e == _T_643 ? $signed(7'shb) : $signed(_GEN_18009); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18011 = 12'h37f == _T_643 ? $signed(7'shc) : $signed(_GEN_18010); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18012 = 12'h380 == _T_643 ? $signed(7'shc) : $signed(_GEN_18011); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18013 = 12'h381 == _T_643 ? $signed(7'shd) : $signed(_GEN_18012); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18014 = 12'h382 == _T_643 ? $signed(7'she) : $signed(_GEN_18013); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18015 = 12'h383 == _T_643 ? $signed(7'shf) : $signed(_GEN_18014); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18016 = 12'h384 == _T_643 ? $signed(7'shf) : $signed(_GEN_18015); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18017 = 12'h385 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18016); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18018 = 12'h386 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18017); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18019 = 12'h387 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18018); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18020 = 12'h388 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18019); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18021 = 12'h389 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18020); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18022 = 12'h38a == _T_643 ? $signed(7'sh14) : $signed(_GEN_18021); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18023 = 12'h38b == _T_643 ? $signed(7'sh14) : $signed(_GEN_18022); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18024 = 12'h38c == _T_643 ? $signed(7'sh15) : $signed(_GEN_18023); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18025 = 12'h38d == _T_643 ? $signed(7'sh16) : $signed(_GEN_18024); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18026 = 12'h38e == _T_643 ? $signed(7'sh16) : $signed(_GEN_18025); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18027 = 12'h38f == _T_643 ? $signed(7'sh17) : $signed(_GEN_18026); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18028 = 12'h390 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18027); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18029 = 12'h391 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18028); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18030 = 12'h392 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18029); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18031 = 12'h393 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18030); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18032 = 12'h394 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18031); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18033 = 12'h395 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18032); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18034 = 12'h396 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18033); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18035 = 12'h397 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18034); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18036 = 12'h398 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_18035); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18037 = 12'h399 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_18036); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18038 = 12'h39a == _T_643 ? $signed(-7'sh1) : $signed(_GEN_18037); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18039 = 12'h39b == _T_643 ? $signed(7'sh0) : $signed(_GEN_18038); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18040 = 12'h39c == _T_643 ? $signed(7'sh0) : $signed(_GEN_18039); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18041 = 12'h39d == _T_643 ? $signed(7'sh1) : $signed(_GEN_18040); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18042 = 12'h39e == _T_643 ? $signed(7'sh2) : $signed(_GEN_18041); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18043 = 12'h39f == _T_643 ? $signed(7'sh3) : $signed(_GEN_18042); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18044 = 12'h3a0 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18043); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18045 = 12'h3a1 == _T_643 ? $signed(7'sh4) : $signed(_GEN_18044); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18046 = 12'h3a2 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18045); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18047 = 12'h3a3 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18046); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18048 = 12'h3a4 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18047); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18049 = 12'h3a5 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18048); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18050 = 12'h3a6 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18049); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18051 = 12'h3a7 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18050); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18052 = 12'h3a8 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18051); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18053 = 12'h3a9 == _T_643 ? $signed(7'sha) : $signed(_GEN_18052); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18054 = 12'h3aa == _T_643 ? $signed(7'sha) : $signed(_GEN_18053); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18055 = 12'h3ab == _T_643 ? $signed(7'shb) : $signed(_GEN_18054); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18056 = 12'h3ac == _T_643 ? $signed(7'shc) : $signed(_GEN_18055); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18057 = 12'h3ad == _T_643 ? $signed(7'shc) : $signed(_GEN_18056); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18058 = 12'h3ae == _T_643 ? $signed(7'shd) : $signed(_GEN_18057); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18059 = 12'h3af == _T_643 ? $signed(7'she) : $signed(_GEN_18058); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18060 = 12'h3b0 == _T_643 ? $signed(7'shf) : $signed(_GEN_18059); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18061 = 12'h3b1 == _T_643 ? $signed(7'shf) : $signed(_GEN_18060); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18062 = 12'h3b2 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18061); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18063 = 12'h3b3 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18062); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18064 = 12'h3b4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18063); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18065 = 12'h3b5 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18064); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18066 = 12'h3b6 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18065); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18067 = 12'h3b7 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18066); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18068 = 12'h3b8 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18067); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18069 = 12'h3b9 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18068); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18070 = 12'h3ba == _T_643 ? $signed(7'sh16) : $signed(_GEN_18069); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18071 = 12'h3bb == _T_643 ? $signed(7'sh16) : $signed(_GEN_18070); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18072 = 12'h3bc == _T_643 ? $signed(7'sh17) : $signed(_GEN_18071); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18073 = 12'h3bd == _T_643 ? $signed(7'sh18) : $signed(_GEN_18072); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18074 = 12'h3be == _T_643 ? $signed(7'sh18) : $signed(_GEN_18073); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18075 = 12'h3bf == _T_643 ? $signed(7'sh19) : $signed(_GEN_18074); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18076 = 12'h3c0 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18075); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18077 = 12'h3c1 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18076); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18078 = 12'h3c2 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18077); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18079 = 12'h3c3 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18078); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18080 = 12'h3c4 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18079); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18081 = 12'h3c5 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18080); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18082 = 12'h3c6 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_18081); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18083 = 12'h3c7 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_18082); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18084 = 12'h3c8 == _T_643 ? $signed(7'sh0) : $signed(_GEN_18083); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18085 = 12'h3c9 == _T_643 ? $signed(7'sh0) : $signed(_GEN_18084); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18086 = 12'h3ca == _T_643 ? $signed(7'sh1) : $signed(_GEN_18085); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18087 = 12'h3cb == _T_643 ? $signed(7'sh2) : $signed(_GEN_18086); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18088 = 12'h3cc == _T_643 ? $signed(7'sh3) : $signed(_GEN_18087); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18089 = 12'h3cd == _T_643 ? $signed(7'sh3) : $signed(_GEN_18088); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18090 = 12'h3ce == _T_643 ? $signed(7'sh4) : $signed(_GEN_18089); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18091 = 12'h3cf == _T_643 ? $signed(7'sh5) : $signed(_GEN_18090); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18092 = 12'h3d0 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18091); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18093 = 12'h3d1 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18092); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18094 = 12'h3d2 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18093); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18095 = 12'h3d3 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18094); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18096 = 12'h3d4 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18095); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18097 = 12'h3d5 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18096); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18098 = 12'h3d6 == _T_643 ? $signed(7'sha) : $signed(_GEN_18097); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18099 = 12'h3d7 == _T_643 ? $signed(7'sha) : $signed(_GEN_18098); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18100 = 12'h3d8 == _T_643 ? $signed(7'shb) : $signed(_GEN_18099); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18101 = 12'h3d9 == _T_643 ? $signed(7'shc) : $signed(_GEN_18100); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18102 = 12'h3da == _T_643 ? $signed(7'shc) : $signed(_GEN_18101); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18103 = 12'h3db == _T_643 ? $signed(7'shd) : $signed(_GEN_18102); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18104 = 12'h3dc == _T_643 ? $signed(7'she) : $signed(_GEN_18103); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18105 = 12'h3dd == _T_643 ? $signed(7'shf) : $signed(_GEN_18104); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18106 = 12'h3de == _T_643 ? $signed(7'shf) : $signed(_GEN_18105); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18107 = 12'h3df == _T_643 ? $signed(7'sh10) : $signed(_GEN_18106); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18108 = 12'h3e0 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18107); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18109 = 12'h3e1 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18108); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18110 = 12'h3e2 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18109); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18111 = 12'h3e3 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18110); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18112 = 12'h3e4 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18111); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18113 = 12'h3e5 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18112); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18114 = 12'h3e6 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18113); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18115 = 12'h3e7 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18114); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18116 = 12'h3e8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18115); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18117 = 12'h3e9 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18116); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18118 = 12'h3ea == _T_643 ? $signed(7'sh18) : $signed(_GEN_18117); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18119 = 12'h3eb == _T_643 ? $signed(7'sh18) : $signed(_GEN_18118); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18120 = 12'h3ec == _T_643 ? $signed(7'sh19) : $signed(_GEN_18119); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18121 = 12'h3ed == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18120); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18122 = 12'h3ee == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18121); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18123 = 12'h3ef == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18122); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18124 = 12'h3f0 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18123); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18125 = 12'h3f1 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18124); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18126 = 12'h3f2 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18125); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18127 = 12'h3f3 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18126); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18128 = 12'h3f4 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_18127); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18129 = 12'h3f5 == _T_643 ? $signed(7'sh0) : $signed(_GEN_18128); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18130 = 12'h3f6 == _T_643 ? $signed(7'sh0) : $signed(_GEN_18129); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18131 = 12'h3f7 == _T_643 ? $signed(7'sh1) : $signed(_GEN_18130); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18132 = 12'h3f8 == _T_643 ? $signed(7'sh2) : $signed(_GEN_18131); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18133 = 12'h3f9 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18132); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18134 = 12'h3fa == _T_643 ? $signed(7'sh3) : $signed(_GEN_18133); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18135 = 12'h3fb == _T_643 ? $signed(7'sh4) : $signed(_GEN_18134); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18136 = 12'h3fc == _T_643 ? $signed(7'sh5) : $signed(_GEN_18135); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18137 = 12'h3fd == _T_643 ? $signed(7'sh5) : $signed(_GEN_18136); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18138 = 12'h3fe == _T_643 ? $signed(7'sh6) : $signed(_GEN_18137); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18139 = 12'h3ff == _T_643 ? $signed(7'sh7) : $signed(_GEN_18138); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18140 = 12'h400 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18139); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18141 = 12'h401 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18140); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18142 = 12'h402 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18141); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18143 = 12'h403 == _T_643 ? $signed(7'sha) : $signed(_GEN_18142); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18144 = 12'h404 == _T_643 ? $signed(7'sha) : $signed(_GEN_18143); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18145 = 12'h405 == _T_643 ? $signed(7'shb) : $signed(_GEN_18144); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18146 = 12'h406 == _T_643 ? $signed(7'shc) : $signed(_GEN_18145); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18147 = 12'h407 == _T_643 ? $signed(7'shc) : $signed(_GEN_18146); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18148 = 12'h408 == _T_643 ? $signed(7'shd) : $signed(_GEN_18147); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18149 = 12'h409 == _T_643 ? $signed(7'she) : $signed(_GEN_18148); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18150 = 12'h40a == _T_643 ? $signed(7'shf) : $signed(_GEN_18149); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18151 = 12'h40b == _T_643 ? $signed(7'shf) : $signed(_GEN_18150); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18152 = 12'h40c == _T_643 ? $signed(7'sh10) : $signed(_GEN_18151); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18153 = 12'h40d == _T_643 ? $signed(7'sh11) : $signed(_GEN_18152); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18154 = 12'h40e == _T_643 ? $signed(7'sh11) : $signed(_GEN_18153); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18155 = 12'h40f == _T_643 ? $signed(7'sh12) : $signed(_GEN_18154); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18156 = 12'h410 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18155); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18157 = 12'h411 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18156); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18158 = 12'h412 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18157); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18159 = 12'h413 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18158); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18160 = 12'h414 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18159); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18161 = 12'h415 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18160); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18162 = 12'h416 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18161); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18163 = 12'h417 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18162); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18164 = 12'h418 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18163); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18165 = 12'h419 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18164); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18166 = 12'h41a == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18165); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18167 = 12'h41b == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18166); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18168 = 12'h41c == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18167); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18169 = 12'h41d == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18168); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18170 = 12'h41e == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18169); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18171 = 12'h41f == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18170); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18172 = 12'h420 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18171); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18173 = 12'h421 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18172); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18174 = 12'h422 == _T_643 ? $signed(7'sh0) : $signed(_GEN_18173); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18175 = 12'h423 == _T_643 ? $signed(7'sh0) : $signed(_GEN_18174); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18176 = 12'h424 == _T_643 ? $signed(7'sh1) : $signed(_GEN_18175); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18177 = 12'h425 == _T_643 ? $signed(7'sh2) : $signed(_GEN_18176); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18178 = 12'h426 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18177); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18179 = 12'h427 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18178); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18180 = 12'h428 == _T_643 ? $signed(7'sh4) : $signed(_GEN_18179); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18181 = 12'h429 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18180); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18182 = 12'h42a == _T_643 ? $signed(7'sh5) : $signed(_GEN_18181); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18183 = 12'h42b == _T_643 ? $signed(7'sh6) : $signed(_GEN_18182); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18184 = 12'h42c == _T_643 ? $signed(7'sh7) : $signed(_GEN_18183); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18185 = 12'h42d == _T_643 ? $signed(7'sh8) : $signed(_GEN_18184); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18186 = 12'h42e == _T_643 ? $signed(7'sh8) : $signed(_GEN_18185); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18187 = 12'h42f == _T_643 ? $signed(7'sh9) : $signed(_GEN_18186); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18188 = 12'h430 == _T_643 ? $signed(7'sha) : $signed(_GEN_18187); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18189 = 12'h431 == _T_643 ? $signed(7'sha) : $signed(_GEN_18188); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18190 = 12'h432 == _T_643 ? $signed(7'shb) : $signed(_GEN_18189); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18191 = 12'h433 == _T_643 ? $signed(7'shc) : $signed(_GEN_18190); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18192 = 12'h434 == _T_643 ? $signed(7'shc) : $signed(_GEN_18191); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18193 = 12'h435 == _T_643 ? $signed(7'shd) : $signed(_GEN_18192); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18194 = 12'h436 == _T_643 ? $signed(7'she) : $signed(_GEN_18193); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18195 = 12'h437 == _T_643 ? $signed(7'shf) : $signed(_GEN_18194); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18196 = 12'h438 == _T_643 ? $signed(7'shf) : $signed(_GEN_18195); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18197 = 12'h439 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18196); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18198 = 12'h43a == _T_643 ? $signed(7'sh11) : $signed(_GEN_18197); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18199 = 12'h43b == _T_643 ? $signed(7'sh11) : $signed(_GEN_18198); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18200 = 12'h43c == _T_643 ? $signed(7'sh12) : $signed(_GEN_18199); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18201 = 12'h43d == _T_643 ? $signed(7'sh13) : $signed(_GEN_18200); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18202 = 12'h43e == _T_643 ? $signed(7'sh14) : $signed(_GEN_18201); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18203 = 12'h43f == _T_643 ? $signed(7'sh14) : $signed(_GEN_18202); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18204 = 12'h440 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18203); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18205 = 12'h441 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18204); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18206 = 12'h442 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18205); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18207 = 12'h443 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18206); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18208 = 12'h444 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18207); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18209 = 12'h445 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18208); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18210 = 12'h446 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18209); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18211 = 12'h447 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18210); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18212 = 12'h448 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18211); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18213 = 12'h449 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18212); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18214 = 12'h44a == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18213); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18215 = 12'h44b == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18214); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18216 = 12'h44c == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18215); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18217 = 12'h44d == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18216); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18218 = 12'h44e == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18217); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18219 = 12'h44f == _T_643 ? $signed(7'sh20) : $signed(_GEN_18218); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18220 = 12'h450 == _T_643 ? $signed(7'sh0) : $signed(_GEN_18219); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18221 = 12'h451 == _T_643 ? $signed(7'sh1) : $signed(_GEN_18220); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18222 = 12'h452 == _T_643 ? $signed(7'sh2) : $signed(_GEN_18221); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18223 = 12'h453 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18222); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18224 = 12'h454 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18223); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18225 = 12'h455 == _T_643 ? $signed(7'sh4) : $signed(_GEN_18224); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18226 = 12'h456 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18225); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18227 = 12'h457 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18226); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18228 = 12'h458 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18227); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18229 = 12'h459 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18228); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18230 = 12'h45a == _T_643 ? $signed(7'sh8) : $signed(_GEN_18229); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18231 = 12'h45b == _T_643 ? $signed(7'sh8) : $signed(_GEN_18230); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18232 = 12'h45c == _T_643 ? $signed(7'sh9) : $signed(_GEN_18231); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18233 = 12'h45d == _T_643 ? $signed(7'sha) : $signed(_GEN_18232); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18234 = 12'h45e == _T_643 ? $signed(7'sha) : $signed(_GEN_18233); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18235 = 12'h45f == _T_643 ? $signed(7'shb) : $signed(_GEN_18234); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18236 = 12'h460 == _T_643 ? $signed(7'shc) : $signed(_GEN_18235); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18237 = 12'h461 == _T_643 ? $signed(7'shc) : $signed(_GEN_18236); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18238 = 12'h462 == _T_643 ? $signed(7'shd) : $signed(_GEN_18237); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18239 = 12'h463 == _T_643 ? $signed(7'she) : $signed(_GEN_18238); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18240 = 12'h464 == _T_643 ? $signed(7'shf) : $signed(_GEN_18239); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18241 = 12'h465 == _T_643 ? $signed(7'shf) : $signed(_GEN_18240); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18242 = 12'h466 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18241); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18243 = 12'h467 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18242); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18244 = 12'h468 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18243); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18245 = 12'h469 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18244); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18246 = 12'h46a == _T_643 ? $signed(7'sh13) : $signed(_GEN_18245); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18247 = 12'h46b == _T_643 ? $signed(7'sh14) : $signed(_GEN_18246); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18248 = 12'h46c == _T_643 ? $signed(7'sh14) : $signed(_GEN_18247); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18249 = 12'h46d == _T_643 ? $signed(7'sh15) : $signed(_GEN_18248); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18250 = 12'h46e == _T_643 ? $signed(7'sh16) : $signed(_GEN_18249); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18251 = 12'h46f == _T_643 ? $signed(7'sh16) : $signed(_GEN_18250); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18252 = 12'h470 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18251); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18253 = 12'h471 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18252); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18254 = 12'h472 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18253); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18255 = 12'h473 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18254); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18256 = 12'h474 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18255); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18257 = 12'h475 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18256); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18258 = 12'h476 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18257); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18259 = 12'h477 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18258); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18260 = 12'h478 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18259); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18261 = 12'h479 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18260); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18262 = 12'h47a == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18261); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18263 = 12'h47b == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18262); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18264 = 12'h47c == _T_643 ? $signed(7'sh20) : $signed(_GEN_18263); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18265 = 12'h47d == _T_643 ? $signed(7'sh20) : $signed(_GEN_18264); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18266 = 12'h47e == _T_643 ? $signed(7'sh1) : $signed(_GEN_18265); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18267 = 12'h47f == _T_643 ? $signed(7'sh2) : $signed(_GEN_18266); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18268 = 12'h480 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18267); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18269 = 12'h481 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18268); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18270 = 12'h482 == _T_643 ? $signed(7'sh4) : $signed(_GEN_18269); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18271 = 12'h483 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18270); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18272 = 12'h484 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18271); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18273 = 12'h485 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18272); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18274 = 12'h486 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18273); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18275 = 12'h487 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18274); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18276 = 12'h488 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18275); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18277 = 12'h489 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18276); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18278 = 12'h48a == _T_643 ? $signed(7'sha) : $signed(_GEN_18277); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18279 = 12'h48b == _T_643 ? $signed(7'sha) : $signed(_GEN_18278); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18280 = 12'h48c == _T_643 ? $signed(7'shb) : $signed(_GEN_18279); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18281 = 12'h48d == _T_643 ? $signed(7'shc) : $signed(_GEN_18280); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18282 = 12'h48e == _T_643 ? $signed(7'shc) : $signed(_GEN_18281); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18283 = 12'h48f == _T_643 ? $signed(7'shd) : $signed(_GEN_18282); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18284 = 12'h490 == _T_643 ? $signed(7'she) : $signed(_GEN_18283); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18285 = 12'h491 == _T_643 ? $signed(7'shf) : $signed(_GEN_18284); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18286 = 12'h492 == _T_643 ? $signed(7'shf) : $signed(_GEN_18285); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18287 = 12'h493 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18286); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18288 = 12'h494 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18287); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18289 = 12'h495 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18288); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18290 = 12'h496 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18289); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18291 = 12'h497 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18290); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18292 = 12'h498 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18291); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18293 = 12'h499 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18292); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18294 = 12'h49a == _T_643 ? $signed(7'sh15) : $signed(_GEN_18293); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18295 = 12'h49b == _T_643 ? $signed(7'sh16) : $signed(_GEN_18294); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18296 = 12'h49c == _T_643 ? $signed(7'sh16) : $signed(_GEN_18295); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18297 = 12'h49d == _T_643 ? $signed(7'sh17) : $signed(_GEN_18296); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18298 = 12'h49e == _T_643 ? $signed(7'sh18) : $signed(_GEN_18297); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18299 = 12'h49f == _T_643 ? $signed(7'sh18) : $signed(_GEN_18298); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18300 = 12'h4a0 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18299); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18301 = 12'h4a1 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18300); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18302 = 12'h4a2 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18301); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18303 = 12'h4a3 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18302); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18304 = 12'h4a4 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18303); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18305 = 12'h4a5 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18304); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18306 = 12'h4a6 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18305); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18307 = 12'h4a7 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18306); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18308 = 12'h4a8 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18307); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18309 = 12'h4a9 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18308); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18310 = 12'h4aa == _T_643 ? $signed(7'sh20) : $signed(_GEN_18309); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18311 = 12'h4ab == _T_643 ? $signed(7'sh21) : $signed(_GEN_18310); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18312 = 12'h4ac == _T_643 ? $signed(7'sh2) : $signed(_GEN_18311); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18313 = 12'h4ad == _T_643 ? $signed(7'sh3) : $signed(_GEN_18312); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18314 = 12'h4ae == _T_643 ? $signed(7'sh3) : $signed(_GEN_18313); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18315 = 12'h4af == _T_643 ? $signed(7'sh4) : $signed(_GEN_18314); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18316 = 12'h4b0 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18315); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18317 = 12'h4b1 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18316); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18318 = 12'h4b2 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18317); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18319 = 12'h4b3 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18318); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18320 = 12'h4b4 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18319); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18321 = 12'h4b5 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18320); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18322 = 12'h4b6 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18321); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18323 = 12'h4b7 == _T_643 ? $signed(7'sha) : $signed(_GEN_18322); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18324 = 12'h4b8 == _T_643 ? $signed(7'sha) : $signed(_GEN_18323); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18325 = 12'h4b9 == _T_643 ? $signed(7'shb) : $signed(_GEN_18324); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18326 = 12'h4ba == _T_643 ? $signed(7'shc) : $signed(_GEN_18325); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18327 = 12'h4bb == _T_643 ? $signed(7'shc) : $signed(_GEN_18326); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18328 = 12'h4bc == _T_643 ? $signed(7'shd) : $signed(_GEN_18327); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18329 = 12'h4bd == _T_643 ? $signed(7'she) : $signed(_GEN_18328); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18330 = 12'h4be == _T_643 ? $signed(7'shf) : $signed(_GEN_18329); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18331 = 12'h4bf == _T_643 ? $signed(7'shf) : $signed(_GEN_18330); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18332 = 12'h4c0 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18331); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18333 = 12'h4c1 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18332); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18334 = 12'h4c2 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18333); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18335 = 12'h4c3 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18334); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18336 = 12'h4c4 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18335); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18337 = 12'h4c5 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18336); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18338 = 12'h4c6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18337); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18339 = 12'h4c7 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18338); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18340 = 12'h4c8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18339); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18341 = 12'h4c9 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18340); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18342 = 12'h4ca == _T_643 ? $signed(7'sh17) : $signed(_GEN_18341); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18343 = 12'h4cb == _T_643 ? $signed(7'sh18) : $signed(_GEN_18342); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18344 = 12'h4cc == _T_643 ? $signed(7'sh18) : $signed(_GEN_18343); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18345 = 12'h4cd == _T_643 ? $signed(7'sh19) : $signed(_GEN_18344); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18346 = 12'h4ce == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18345); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18347 = 12'h4cf == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18346); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18348 = 12'h4d0 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18347); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18349 = 12'h4d1 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18348); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18350 = 12'h4d2 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18349); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18351 = 12'h4d3 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18350); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18352 = 12'h4d4 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18351); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18353 = 12'h4d5 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18352); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18354 = 12'h4d6 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18353); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18355 = 12'h4d7 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18354); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18356 = 12'h4d8 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18355); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18357 = 12'h4d9 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18356); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18358 = 12'h4da == _T_643 ? $signed(7'sh3) : $signed(_GEN_18357); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18359 = 12'h4db == _T_643 ? $signed(7'sh3) : $signed(_GEN_18358); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18360 = 12'h4dc == _T_643 ? $signed(7'sh4) : $signed(_GEN_18359); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18361 = 12'h4dd == _T_643 ? $signed(7'sh5) : $signed(_GEN_18360); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18362 = 12'h4de == _T_643 ? $signed(7'sh5) : $signed(_GEN_18361); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18363 = 12'h4df == _T_643 ? $signed(7'sh6) : $signed(_GEN_18362); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18364 = 12'h4e0 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18363); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18365 = 12'h4e1 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18364); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18366 = 12'h4e2 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18365); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18367 = 12'h4e3 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18366); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18368 = 12'h4e4 == _T_643 ? $signed(7'sha) : $signed(_GEN_18367); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18369 = 12'h4e5 == _T_643 ? $signed(7'sha) : $signed(_GEN_18368); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18370 = 12'h4e6 == _T_643 ? $signed(7'shb) : $signed(_GEN_18369); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18371 = 12'h4e7 == _T_643 ? $signed(7'shc) : $signed(_GEN_18370); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18372 = 12'h4e8 == _T_643 ? $signed(7'shc) : $signed(_GEN_18371); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18373 = 12'h4e9 == _T_643 ? $signed(7'shd) : $signed(_GEN_18372); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18374 = 12'h4ea == _T_643 ? $signed(7'she) : $signed(_GEN_18373); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18375 = 12'h4eb == _T_643 ? $signed(7'shf) : $signed(_GEN_18374); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18376 = 12'h4ec == _T_643 ? $signed(7'shf) : $signed(_GEN_18375); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18377 = 12'h4ed == _T_643 ? $signed(7'sh10) : $signed(_GEN_18376); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18378 = 12'h4ee == _T_643 ? $signed(7'sh11) : $signed(_GEN_18377); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18379 = 12'h4ef == _T_643 ? $signed(7'sh11) : $signed(_GEN_18378); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18380 = 12'h4f0 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18379); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18381 = 12'h4f1 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18380); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18382 = 12'h4f2 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18381); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18383 = 12'h4f3 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18382); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18384 = 12'h4f4 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18383); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18385 = 12'h4f5 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18384); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18386 = 12'h4f6 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18385); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18387 = 12'h4f7 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18386); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18388 = 12'h4f8 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18387); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18389 = 12'h4f9 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18388); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18390 = 12'h4fa == _T_643 ? $signed(7'sh19) : $signed(_GEN_18389); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18391 = 12'h4fb == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18390); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18392 = 12'h4fc == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18391); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18393 = 12'h4fd == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18392); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18394 = 12'h4fe == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18393); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18395 = 12'h4ff == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18394); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18396 = 12'h500 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18395); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18397 = 12'h501 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18396); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18398 = 12'h502 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18397); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18399 = 12'h503 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18398); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18400 = 12'h504 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18399); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18401 = 12'h505 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18400); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18402 = 12'h506 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18401); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18403 = 12'h507 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18402); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18404 = 12'h508 == _T_643 ? $signed(7'sh3) : $signed(_GEN_18403); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18405 = 12'h509 == _T_643 ? $signed(7'sh4) : $signed(_GEN_18404); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18406 = 12'h50a == _T_643 ? $signed(7'sh5) : $signed(_GEN_18405); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18407 = 12'h50b == _T_643 ? $signed(7'sh5) : $signed(_GEN_18406); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18408 = 12'h50c == _T_643 ? $signed(7'sh6) : $signed(_GEN_18407); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18409 = 12'h50d == _T_643 ? $signed(7'sh7) : $signed(_GEN_18408); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18410 = 12'h50e == _T_643 ? $signed(7'sh8) : $signed(_GEN_18409); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18411 = 12'h50f == _T_643 ? $signed(7'sh8) : $signed(_GEN_18410); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18412 = 12'h510 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18411); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18413 = 12'h511 == _T_643 ? $signed(7'sha) : $signed(_GEN_18412); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18414 = 12'h512 == _T_643 ? $signed(7'sha) : $signed(_GEN_18413); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18415 = 12'h513 == _T_643 ? $signed(7'shb) : $signed(_GEN_18414); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18416 = 12'h514 == _T_643 ? $signed(7'shc) : $signed(_GEN_18415); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18417 = 12'h515 == _T_643 ? $signed(7'shc) : $signed(_GEN_18416); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18418 = 12'h516 == _T_643 ? $signed(7'shd) : $signed(_GEN_18417); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18419 = 12'h517 == _T_643 ? $signed(7'she) : $signed(_GEN_18418); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18420 = 12'h518 == _T_643 ? $signed(7'shf) : $signed(_GEN_18419); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18421 = 12'h519 == _T_643 ? $signed(7'shf) : $signed(_GEN_18420); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18422 = 12'h51a == _T_643 ? $signed(7'sh10) : $signed(_GEN_18421); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18423 = 12'h51b == _T_643 ? $signed(7'sh11) : $signed(_GEN_18422); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18424 = 12'h51c == _T_643 ? $signed(7'sh11) : $signed(_GEN_18423); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18425 = 12'h51d == _T_643 ? $signed(7'sh12) : $signed(_GEN_18424); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18426 = 12'h51e == _T_643 ? $signed(7'sh13) : $signed(_GEN_18425); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18427 = 12'h51f == _T_643 ? $signed(7'sh14) : $signed(_GEN_18426); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18428 = 12'h520 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18427); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18429 = 12'h521 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18428); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18430 = 12'h522 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18429); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18431 = 12'h523 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18430); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18432 = 12'h524 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18431); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18433 = 12'h525 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18432); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18434 = 12'h526 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18433); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18435 = 12'h527 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18434); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18436 = 12'h528 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18435); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18437 = 12'h529 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18436); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18438 = 12'h52a == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18437); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18439 = 12'h52b == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18438); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18440 = 12'h52c == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18439); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18441 = 12'h52d == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18440); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18442 = 12'h52e == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18441); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18443 = 12'h52f == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18442); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18444 = 12'h530 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18443); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18445 = 12'h531 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18444); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18446 = 12'h532 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18445); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18447 = 12'h533 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18446); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18448 = 12'h534 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18447); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18449 = 12'h535 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18448); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18450 = 12'h536 == _T_643 ? $signed(7'sh4) : $signed(_GEN_18449); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18451 = 12'h537 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18450); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18452 = 12'h538 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18451); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18453 = 12'h539 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18452); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18454 = 12'h53a == _T_643 ? $signed(7'sh7) : $signed(_GEN_18453); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18455 = 12'h53b == _T_643 ? $signed(7'sh8) : $signed(_GEN_18454); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18456 = 12'h53c == _T_643 ? $signed(7'sh8) : $signed(_GEN_18455); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18457 = 12'h53d == _T_643 ? $signed(7'sh9) : $signed(_GEN_18456); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18458 = 12'h53e == _T_643 ? $signed(7'sha) : $signed(_GEN_18457); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18459 = 12'h53f == _T_643 ? $signed(7'sha) : $signed(_GEN_18458); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18460 = 12'h540 == _T_643 ? $signed(7'shb) : $signed(_GEN_18459); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18461 = 12'h541 == _T_643 ? $signed(7'shc) : $signed(_GEN_18460); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18462 = 12'h542 == _T_643 ? $signed(7'shc) : $signed(_GEN_18461); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18463 = 12'h543 == _T_643 ? $signed(7'shd) : $signed(_GEN_18462); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18464 = 12'h544 == _T_643 ? $signed(7'she) : $signed(_GEN_18463); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18465 = 12'h545 == _T_643 ? $signed(7'shf) : $signed(_GEN_18464); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18466 = 12'h546 == _T_643 ? $signed(7'shf) : $signed(_GEN_18465); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18467 = 12'h547 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18466); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18468 = 12'h548 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18467); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18469 = 12'h549 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18468); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18470 = 12'h54a == _T_643 ? $signed(7'sh12) : $signed(_GEN_18469); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18471 = 12'h54b == _T_643 ? $signed(7'sh13) : $signed(_GEN_18470); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18472 = 12'h54c == _T_643 ? $signed(7'sh14) : $signed(_GEN_18471); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18473 = 12'h54d == _T_643 ? $signed(7'sh14) : $signed(_GEN_18472); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18474 = 12'h54e == _T_643 ? $signed(7'sh15) : $signed(_GEN_18473); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18475 = 12'h54f == _T_643 ? $signed(7'sh16) : $signed(_GEN_18474); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18476 = 12'h550 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18475); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18477 = 12'h551 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18476); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18478 = 12'h552 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18477); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18479 = 12'h553 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18478); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18480 = 12'h554 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18479); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18481 = 12'h555 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18480); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18482 = 12'h556 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18481); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18483 = 12'h557 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18482); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18484 = 12'h558 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18483); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18485 = 12'h559 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18484); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18486 = 12'h55a == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18485); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18487 = 12'h55b == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18486); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18488 = 12'h55c == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18487); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18489 = 12'h55d == _T_643 ? $signed(7'sh20) : $signed(_GEN_18488); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18490 = 12'h55e == _T_643 ? $signed(7'sh20) : $signed(_GEN_18489); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18491 = 12'h55f == _T_643 ? $signed(7'sh21) : $signed(_GEN_18490); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18492 = 12'h560 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18491); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18493 = 12'h561 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18492); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18494 = 12'h562 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18493); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18495 = 12'h563 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18494); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18496 = 12'h564 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18495); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18497 = 12'h565 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18496); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18498 = 12'h566 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18497); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18499 = 12'h567 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18498); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18500 = 12'h568 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18499); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18501 = 12'h569 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18500); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18502 = 12'h56a == _T_643 ? $signed(7'sh9) : $signed(_GEN_18501); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18503 = 12'h56b == _T_643 ? $signed(7'sha) : $signed(_GEN_18502); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18504 = 12'h56c == _T_643 ? $signed(7'sha) : $signed(_GEN_18503); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18505 = 12'h56d == _T_643 ? $signed(7'shb) : $signed(_GEN_18504); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18506 = 12'h56e == _T_643 ? $signed(7'shc) : $signed(_GEN_18505); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18507 = 12'h56f == _T_643 ? $signed(7'shc) : $signed(_GEN_18506); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18508 = 12'h570 == _T_643 ? $signed(7'shd) : $signed(_GEN_18507); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18509 = 12'h571 == _T_643 ? $signed(7'she) : $signed(_GEN_18508); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18510 = 12'h572 == _T_643 ? $signed(7'shf) : $signed(_GEN_18509); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18511 = 12'h573 == _T_643 ? $signed(7'shf) : $signed(_GEN_18510); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18512 = 12'h574 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18511); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18513 = 12'h575 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18512); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18514 = 12'h576 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18513); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18515 = 12'h577 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18514); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18516 = 12'h578 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18515); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18517 = 12'h579 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18516); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18518 = 12'h57a == _T_643 ? $signed(7'sh14) : $signed(_GEN_18517); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18519 = 12'h57b == _T_643 ? $signed(7'sh15) : $signed(_GEN_18518); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18520 = 12'h57c == _T_643 ? $signed(7'sh16) : $signed(_GEN_18519); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18521 = 12'h57d == _T_643 ? $signed(7'sh16) : $signed(_GEN_18520); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18522 = 12'h57e == _T_643 ? $signed(7'sh17) : $signed(_GEN_18521); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18523 = 12'h57f == _T_643 ? $signed(7'sh18) : $signed(_GEN_18522); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18524 = 12'h580 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18523); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18525 = 12'h581 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18524); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18526 = 12'h582 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18525); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18527 = 12'h583 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18526); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18528 = 12'h584 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18527); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18529 = 12'h585 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18528); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18530 = 12'h586 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18529); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18531 = 12'h587 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18530); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18532 = 12'h588 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18531); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18533 = 12'h589 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18532); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18534 = 12'h58a == _T_643 ? $signed(7'sh20) : $signed(_GEN_18533); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18535 = 12'h58b == _T_643 ? $signed(7'sh20) : $signed(_GEN_18534); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18536 = 12'h58c == _T_643 ? $signed(7'sh21) : $signed(_GEN_18535); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18537 = 12'h58d == _T_643 ? $signed(7'sh22) : $signed(_GEN_18536); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18538 = 12'h58e == _T_643 ? $signed(7'sh22) : $signed(_GEN_18537); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18539 = 12'h58f == _T_643 ? $signed(7'sh23) : $signed(_GEN_18538); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18540 = 12'h590 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18539); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18541 = 12'h591 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18540); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18542 = 12'h592 == _T_643 ? $signed(7'sh5) : $signed(_GEN_18541); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18543 = 12'h593 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18542); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18544 = 12'h594 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18543); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18545 = 12'h595 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18544); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18546 = 12'h596 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18545); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18547 = 12'h597 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18546); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18548 = 12'h598 == _T_643 ? $signed(7'sha) : $signed(_GEN_18547); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18549 = 12'h599 == _T_643 ? $signed(7'sha) : $signed(_GEN_18548); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18550 = 12'h59a == _T_643 ? $signed(7'shb) : $signed(_GEN_18549); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18551 = 12'h59b == _T_643 ? $signed(7'shc) : $signed(_GEN_18550); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18552 = 12'h59c == _T_643 ? $signed(7'shc) : $signed(_GEN_18551); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18553 = 12'h59d == _T_643 ? $signed(7'shd) : $signed(_GEN_18552); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18554 = 12'h59e == _T_643 ? $signed(7'she) : $signed(_GEN_18553); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18555 = 12'h59f == _T_643 ? $signed(7'shf) : $signed(_GEN_18554); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18556 = 12'h5a0 == _T_643 ? $signed(7'shf) : $signed(_GEN_18555); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18557 = 12'h5a1 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18556); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18558 = 12'h5a2 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18557); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18559 = 12'h5a3 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18558); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18560 = 12'h5a4 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18559); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18561 = 12'h5a5 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18560); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18562 = 12'h5a6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18561); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18563 = 12'h5a7 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18562); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18564 = 12'h5a8 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18563); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18565 = 12'h5a9 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18564); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18566 = 12'h5aa == _T_643 ? $signed(7'sh16) : $signed(_GEN_18565); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18567 = 12'h5ab == _T_643 ? $signed(7'sh17) : $signed(_GEN_18566); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18568 = 12'h5ac == _T_643 ? $signed(7'sh18) : $signed(_GEN_18567); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18569 = 12'h5ad == _T_643 ? $signed(7'sh18) : $signed(_GEN_18568); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18570 = 12'h5ae == _T_643 ? $signed(7'sh19) : $signed(_GEN_18569); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18571 = 12'h5af == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18570); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18572 = 12'h5b0 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18571); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18573 = 12'h5b1 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18572); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18574 = 12'h5b2 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18573); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18575 = 12'h5b3 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18574); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18576 = 12'h5b4 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18575); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18577 = 12'h5b5 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18576); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18578 = 12'h5b6 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18577); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18579 = 12'h5b7 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18578); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18580 = 12'h5b8 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18579); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18581 = 12'h5b9 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18580); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18582 = 12'h5ba == _T_643 ? $signed(7'sh22) : $signed(_GEN_18581); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18583 = 12'h5bb == _T_643 ? $signed(7'sh22) : $signed(_GEN_18582); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18584 = 12'h5bc == _T_643 ? $signed(7'sh23) : $signed(_GEN_18583); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18585 = 12'h5bd == _T_643 ? $signed(7'sh24) : $signed(_GEN_18584); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18586 = 12'h5be == _T_643 ? $signed(7'sh25) : $signed(_GEN_18585); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18587 = 12'h5bf == _T_643 ? $signed(7'sh25) : $signed(_GEN_18586); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18588 = 12'h5c0 == _T_643 ? $signed(7'sh6) : $signed(_GEN_18587); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18589 = 12'h5c1 == _T_643 ? $signed(7'sh7) : $signed(_GEN_18588); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18590 = 12'h5c2 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18589); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18591 = 12'h5c3 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18590); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18592 = 12'h5c4 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18591); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18593 = 12'h5c5 == _T_643 ? $signed(7'sha) : $signed(_GEN_18592); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18594 = 12'h5c6 == _T_643 ? $signed(7'sha) : $signed(_GEN_18593); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18595 = 12'h5c7 == _T_643 ? $signed(7'shb) : $signed(_GEN_18594); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18596 = 12'h5c8 == _T_643 ? $signed(7'shc) : $signed(_GEN_18595); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18597 = 12'h5c9 == _T_643 ? $signed(7'shc) : $signed(_GEN_18596); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18598 = 12'h5ca == _T_643 ? $signed(7'shd) : $signed(_GEN_18597); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18599 = 12'h5cb == _T_643 ? $signed(7'she) : $signed(_GEN_18598); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18600 = 12'h5cc == _T_643 ? $signed(7'shf) : $signed(_GEN_18599); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18601 = 12'h5cd == _T_643 ? $signed(7'shf) : $signed(_GEN_18600); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18602 = 12'h5ce == _T_643 ? $signed(7'sh10) : $signed(_GEN_18601); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18603 = 12'h5cf == _T_643 ? $signed(7'sh11) : $signed(_GEN_18602); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18604 = 12'h5d0 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18603); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18605 = 12'h5d1 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18604); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18606 = 12'h5d2 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18605); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18607 = 12'h5d3 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18606); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18608 = 12'h5d4 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18607); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18609 = 12'h5d5 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18608); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18610 = 12'h5d6 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18609); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18611 = 12'h5d7 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18610); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18612 = 12'h5d8 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18611); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18613 = 12'h5d9 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18612); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18614 = 12'h5da == _T_643 ? $signed(7'sh18) : $signed(_GEN_18613); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18615 = 12'h5db == _T_643 ? $signed(7'sh19) : $signed(_GEN_18614); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18616 = 12'h5dc == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18615); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18617 = 12'h5dd == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18616); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18618 = 12'h5de == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18617); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18619 = 12'h5df == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18618); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18620 = 12'h5e0 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18619); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18621 = 12'h5e1 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18620); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18622 = 12'h5e2 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18621); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18623 = 12'h5e3 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18622); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18624 = 12'h5e4 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18623); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18625 = 12'h5e5 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18624); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18626 = 12'h5e6 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18625); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18627 = 12'h5e7 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18626); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18628 = 12'h5e8 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18627); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18629 = 12'h5e9 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18628); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18630 = 12'h5ea == _T_643 ? $signed(7'sh24) : $signed(_GEN_18629); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18631 = 12'h5eb == _T_643 ? $signed(7'sh25) : $signed(_GEN_18630); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18632 = 12'h5ec == _T_643 ? $signed(7'sh25) : $signed(_GEN_18631); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18633 = 12'h5ed == _T_643 ? $signed(7'sh26) : $signed(_GEN_18632); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18634 = 12'h5ee == _T_643 ? $signed(7'sh7) : $signed(_GEN_18633); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18635 = 12'h5ef == _T_643 ? $signed(7'sh8) : $signed(_GEN_18634); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18636 = 12'h5f0 == _T_643 ? $signed(7'sh8) : $signed(_GEN_18635); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18637 = 12'h5f1 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18636); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18638 = 12'h5f2 == _T_643 ? $signed(7'sha) : $signed(_GEN_18637); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18639 = 12'h5f3 == _T_643 ? $signed(7'sha) : $signed(_GEN_18638); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18640 = 12'h5f4 == _T_643 ? $signed(7'shb) : $signed(_GEN_18639); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18641 = 12'h5f5 == _T_643 ? $signed(7'shc) : $signed(_GEN_18640); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18642 = 12'h5f6 == _T_643 ? $signed(7'shc) : $signed(_GEN_18641); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18643 = 12'h5f7 == _T_643 ? $signed(7'shd) : $signed(_GEN_18642); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18644 = 12'h5f8 == _T_643 ? $signed(7'she) : $signed(_GEN_18643); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18645 = 12'h5f9 == _T_643 ? $signed(7'shf) : $signed(_GEN_18644); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18646 = 12'h5fa == _T_643 ? $signed(7'shf) : $signed(_GEN_18645); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18647 = 12'h5fb == _T_643 ? $signed(7'sh10) : $signed(_GEN_18646); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18648 = 12'h5fc == _T_643 ? $signed(7'sh11) : $signed(_GEN_18647); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18649 = 12'h5fd == _T_643 ? $signed(7'sh11) : $signed(_GEN_18648); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18650 = 12'h5fe == _T_643 ? $signed(7'sh12) : $signed(_GEN_18649); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18651 = 12'h5ff == _T_643 ? $signed(7'sh13) : $signed(_GEN_18650); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18652 = 12'h600 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18651); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18653 = 12'h601 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18652); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18654 = 12'h602 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18653); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18655 = 12'h603 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18654); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18656 = 12'h604 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18655); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18657 = 12'h605 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18656); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18658 = 12'h606 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18657); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18659 = 12'h607 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18658); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18660 = 12'h608 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18659); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18661 = 12'h609 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18660); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18662 = 12'h60a == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18661); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18663 = 12'h60b == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18662); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18664 = 12'h60c == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18663); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18665 = 12'h60d == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18664); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18666 = 12'h60e == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18665); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18667 = 12'h60f == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18666); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18668 = 12'h610 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18667); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18669 = 12'h611 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18668); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18670 = 12'h612 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18669); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18671 = 12'h613 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18670); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18672 = 12'h614 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18671); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18673 = 12'h615 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18672); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18674 = 12'h616 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18673); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18675 = 12'h617 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18674); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18676 = 12'h618 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18675); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18677 = 12'h619 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18676); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18678 = 12'h61a == _T_643 ? $signed(7'sh26) : $signed(_GEN_18677); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18679 = 12'h61b == _T_643 ? $signed(7'sh27) : $signed(_GEN_18678); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18680 = 12'h61c == _T_643 ? $signed(7'sh8) : $signed(_GEN_18679); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18681 = 12'h61d == _T_643 ? $signed(7'sh8) : $signed(_GEN_18680); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18682 = 12'h61e == _T_643 ? $signed(7'sh9) : $signed(_GEN_18681); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18683 = 12'h61f == _T_643 ? $signed(7'sha) : $signed(_GEN_18682); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18684 = 12'h620 == _T_643 ? $signed(7'sha) : $signed(_GEN_18683); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18685 = 12'h621 == _T_643 ? $signed(7'shb) : $signed(_GEN_18684); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18686 = 12'h622 == _T_643 ? $signed(7'shc) : $signed(_GEN_18685); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18687 = 12'h623 == _T_643 ? $signed(7'shc) : $signed(_GEN_18686); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18688 = 12'h624 == _T_643 ? $signed(7'shd) : $signed(_GEN_18687); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18689 = 12'h625 == _T_643 ? $signed(7'she) : $signed(_GEN_18688); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18690 = 12'h626 == _T_643 ? $signed(7'shf) : $signed(_GEN_18689); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18691 = 12'h627 == _T_643 ? $signed(7'shf) : $signed(_GEN_18690); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18692 = 12'h628 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18691); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18693 = 12'h629 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18692); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18694 = 12'h62a == _T_643 ? $signed(7'sh11) : $signed(_GEN_18693); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18695 = 12'h62b == _T_643 ? $signed(7'sh12) : $signed(_GEN_18694); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18696 = 12'h62c == _T_643 ? $signed(7'sh13) : $signed(_GEN_18695); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18697 = 12'h62d == _T_643 ? $signed(7'sh14) : $signed(_GEN_18696); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18698 = 12'h62e == _T_643 ? $signed(7'sh14) : $signed(_GEN_18697); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18699 = 12'h62f == _T_643 ? $signed(7'sh15) : $signed(_GEN_18698); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18700 = 12'h630 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18699); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18701 = 12'h631 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18700); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18702 = 12'h632 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18701); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18703 = 12'h633 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18702); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18704 = 12'h634 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18703); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18705 = 12'h635 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18704); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18706 = 12'h636 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18705); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18707 = 12'h637 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18706); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18708 = 12'h638 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18707); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18709 = 12'h639 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18708); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18710 = 12'h63a == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18709); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18711 = 12'h63b == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18710); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18712 = 12'h63c == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18711); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18713 = 12'h63d == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18712); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18714 = 12'h63e == _T_643 ? $signed(7'sh20) : $signed(_GEN_18713); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18715 = 12'h63f == _T_643 ? $signed(7'sh20) : $signed(_GEN_18714); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18716 = 12'h640 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18715); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18717 = 12'h641 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18716); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18718 = 12'h642 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18717); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18719 = 12'h643 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18718); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18720 = 12'h644 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18719); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18721 = 12'h645 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18720); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18722 = 12'h646 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18721); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18723 = 12'h647 == _T_643 ? $signed(7'sh26) : $signed(_GEN_18722); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18724 = 12'h648 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18723); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18725 = 12'h649 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18724); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18726 = 12'h64a == _T_643 ? $signed(7'sh8) : $signed(_GEN_18725); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18727 = 12'h64b == _T_643 ? $signed(7'sh9) : $signed(_GEN_18726); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18728 = 12'h64c == _T_643 ? $signed(7'sha) : $signed(_GEN_18727); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18729 = 12'h64d == _T_643 ? $signed(7'sha) : $signed(_GEN_18728); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18730 = 12'h64e == _T_643 ? $signed(7'shb) : $signed(_GEN_18729); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18731 = 12'h64f == _T_643 ? $signed(7'shc) : $signed(_GEN_18730); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18732 = 12'h650 == _T_643 ? $signed(7'shc) : $signed(_GEN_18731); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18733 = 12'h651 == _T_643 ? $signed(7'shd) : $signed(_GEN_18732); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18734 = 12'h652 == _T_643 ? $signed(7'she) : $signed(_GEN_18733); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18735 = 12'h653 == _T_643 ? $signed(7'shf) : $signed(_GEN_18734); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18736 = 12'h654 == _T_643 ? $signed(7'shf) : $signed(_GEN_18735); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18737 = 12'h655 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18736); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18738 = 12'h656 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18737); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18739 = 12'h657 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18738); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18740 = 12'h658 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18739); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18741 = 12'h659 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18740); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18742 = 12'h65a == _T_643 ? $signed(7'sh14) : $signed(_GEN_18741); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18743 = 12'h65b == _T_643 ? $signed(7'sh14) : $signed(_GEN_18742); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18744 = 12'h65c == _T_643 ? $signed(7'sh15) : $signed(_GEN_18743); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18745 = 12'h65d == _T_643 ? $signed(7'sh16) : $signed(_GEN_18744); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18746 = 12'h65e == _T_643 ? $signed(7'sh16) : $signed(_GEN_18745); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18747 = 12'h65f == _T_643 ? $signed(7'sh17) : $signed(_GEN_18746); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18748 = 12'h660 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18747); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18749 = 12'h661 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18748); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18750 = 12'h662 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18749); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18751 = 12'h663 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18750); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18752 = 12'h664 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18751); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18753 = 12'h665 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18752); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18754 = 12'h666 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18753); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18755 = 12'h667 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18754); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18756 = 12'h668 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18755); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18757 = 12'h669 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18756); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18758 = 12'h66a == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18757); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18759 = 12'h66b == _T_643 ? $signed(7'sh20) : $signed(_GEN_18758); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18760 = 12'h66c == _T_643 ? $signed(7'sh20) : $signed(_GEN_18759); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18761 = 12'h66d == _T_643 ? $signed(7'sh21) : $signed(_GEN_18760); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18762 = 12'h66e == _T_643 ? $signed(7'sh22) : $signed(_GEN_18761); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18763 = 12'h66f == _T_643 ? $signed(7'sh22) : $signed(_GEN_18762); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18764 = 12'h670 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18763); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18765 = 12'h671 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18764); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18766 = 12'h672 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18765); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18767 = 12'h673 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18766); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18768 = 12'h674 == _T_643 ? $signed(7'sh26) : $signed(_GEN_18767); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18769 = 12'h675 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18768); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18770 = 12'h676 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18769); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18771 = 12'h677 == _T_643 ? $signed(7'sh28) : $signed(_GEN_18770); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18772 = 12'h678 == _T_643 ? $signed(7'sh9) : $signed(_GEN_18771); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18773 = 12'h679 == _T_643 ? $signed(7'sha) : $signed(_GEN_18772); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18774 = 12'h67a == _T_643 ? $signed(7'sha) : $signed(_GEN_18773); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18775 = 12'h67b == _T_643 ? $signed(7'shb) : $signed(_GEN_18774); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18776 = 12'h67c == _T_643 ? $signed(7'shc) : $signed(_GEN_18775); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18777 = 12'h67d == _T_643 ? $signed(7'shc) : $signed(_GEN_18776); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18778 = 12'h67e == _T_643 ? $signed(7'shd) : $signed(_GEN_18777); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18779 = 12'h67f == _T_643 ? $signed(7'she) : $signed(_GEN_18778); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18780 = 12'h680 == _T_643 ? $signed(7'shf) : $signed(_GEN_18779); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18781 = 12'h681 == _T_643 ? $signed(7'shf) : $signed(_GEN_18780); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18782 = 12'h682 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18781); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18783 = 12'h683 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18782); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18784 = 12'h684 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18783); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18785 = 12'h685 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18784); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18786 = 12'h686 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18785); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18787 = 12'h687 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18786); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18788 = 12'h688 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18787); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18789 = 12'h689 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18788); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18790 = 12'h68a == _T_643 ? $signed(7'sh16) : $signed(_GEN_18789); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18791 = 12'h68b == _T_643 ? $signed(7'sh16) : $signed(_GEN_18790); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18792 = 12'h68c == _T_643 ? $signed(7'sh17) : $signed(_GEN_18791); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18793 = 12'h68d == _T_643 ? $signed(7'sh18) : $signed(_GEN_18792); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18794 = 12'h68e == _T_643 ? $signed(7'sh18) : $signed(_GEN_18793); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18795 = 12'h68f == _T_643 ? $signed(7'sh19) : $signed(_GEN_18794); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18796 = 12'h690 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18795); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18797 = 12'h691 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18796); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18798 = 12'h692 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18797); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18799 = 12'h693 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18798); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18800 = 12'h694 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18799); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18801 = 12'h695 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18800); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18802 = 12'h696 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18801); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18803 = 12'h697 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18802); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18804 = 12'h698 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18803); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18805 = 12'h699 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18804); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18806 = 12'h69a == _T_643 ? $signed(7'sh21) : $signed(_GEN_18805); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18807 = 12'h69b == _T_643 ? $signed(7'sh22) : $signed(_GEN_18806); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18808 = 12'h69c == _T_643 ? $signed(7'sh22) : $signed(_GEN_18807); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18809 = 12'h69d == _T_643 ? $signed(7'sh23) : $signed(_GEN_18808); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18810 = 12'h69e == _T_643 ? $signed(7'sh24) : $signed(_GEN_18809); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18811 = 12'h69f == _T_643 ? $signed(7'sh25) : $signed(_GEN_18810); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18812 = 12'h6a0 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18811); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18813 = 12'h6a1 == _T_643 ? $signed(7'sh26) : $signed(_GEN_18812); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18814 = 12'h6a2 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18813); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18815 = 12'h6a3 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18814); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18816 = 12'h6a4 == _T_643 ? $signed(7'sh28) : $signed(_GEN_18815); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18817 = 12'h6a5 == _T_643 ? $signed(7'sh29) : $signed(_GEN_18816); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18818 = 12'h6a6 == _T_643 ? $signed(7'sha) : $signed(_GEN_18817); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18819 = 12'h6a7 == _T_643 ? $signed(7'sha) : $signed(_GEN_18818); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18820 = 12'h6a8 == _T_643 ? $signed(7'shb) : $signed(_GEN_18819); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18821 = 12'h6a9 == _T_643 ? $signed(7'shc) : $signed(_GEN_18820); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18822 = 12'h6aa == _T_643 ? $signed(7'shc) : $signed(_GEN_18821); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18823 = 12'h6ab == _T_643 ? $signed(7'shd) : $signed(_GEN_18822); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18824 = 12'h6ac == _T_643 ? $signed(7'she) : $signed(_GEN_18823); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18825 = 12'h6ad == _T_643 ? $signed(7'shf) : $signed(_GEN_18824); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18826 = 12'h6ae == _T_643 ? $signed(7'shf) : $signed(_GEN_18825); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18827 = 12'h6af == _T_643 ? $signed(7'sh10) : $signed(_GEN_18826); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18828 = 12'h6b0 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18827); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18829 = 12'h6b1 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18828); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18830 = 12'h6b2 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18829); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18831 = 12'h6b3 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18830); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18832 = 12'h6b4 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18831); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18833 = 12'h6b5 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18832); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18834 = 12'h6b6 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18833); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18835 = 12'h6b7 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18834); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18836 = 12'h6b8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18835); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18837 = 12'h6b9 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18836); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18838 = 12'h6ba == _T_643 ? $signed(7'sh18) : $signed(_GEN_18837); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18839 = 12'h6bb == _T_643 ? $signed(7'sh18) : $signed(_GEN_18838); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18840 = 12'h6bc == _T_643 ? $signed(7'sh19) : $signed(_GEN_18839); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18841 = 12'h6bd == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18840); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18842 = 12'h6be == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18841); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18843 = 12'h6bf == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18842); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18844 = 12'h6c0 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18843); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18845 = 12'h6c1 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18844); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18846 = 12'h6c2 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18845); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18847 = 12'h6c3 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18846); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18848 = 12'h6c4 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18847); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18849 = 12'h6c5 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18848); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18850 = 12'h6c6 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18849); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18851 = 12'h6c7 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18850); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18852 = 12'h6c8 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18851); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18853 = 12'h6c9 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18852); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18854 = 12'h6ca == _T_643 ? $signed(7'sh23) : $signed(_GEN_18853); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18855 = 12'h6cb == _T_643 ? $signed(7'sh24) : $signed(_GEN_18854); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18856 = 12'h6cc == _T_643 ? $signed(7'sh25) : $signed(_GEN_18855); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18857 = 12'h6cd == _T_643 ? $signed(7'sh25) : $signed(_GEN_18856); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18858 = 12'h6ce == _T_643 ? $signed(7'sh26) : $signed(_GEN_18857); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18859 = 12'h6cf == _T_643 ? $signed(7'sh27) : $signed(_GEN_18858); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18860 = 12'h6d0 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18859); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18861 = 12'h6d1 == _T_643 ? $signed(7'sh28) : $signed(_GEN_18860); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18862 = 12'h6d2 == _T_643 ? $signed(7'sh29) : $signed(_GEN_18861); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18863 = 12'h6d3 == _T_643 ? $signed(7'sh29) : $signed(_GEN_18862); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18864 = 12'h6d4 == _T_643 ? $signed(7'sha) : $signed(_GEN_18863); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18865 = 12'h6d5 == _T_643 ? $signed(7'shb) : $signed(_GEN_18864); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18866 = 12'h6d6 == _T_643 ? $signed(7'shc) : $signed(_GEN_18865); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18867 = 12'h6d7 == _T_643 ? $signed(7'shc) : $signed(_GEN_18866); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18868 = 12'h6d8 == _T_643 ? $signed(7'shd) : $signed(_GEN_18867); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18869 = 12'h6d9 == _T_643 ? $signed(7'she) : $signed(_GEN_18868); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18870 = 12'h6da == _T_643 ? $signed(7'shf) : $signed(_GEN_18869); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18871 = 12'h6db == _T_643 ? $signed(7'shf) : $signed(_GEN_18870); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18872 = 12'h6dc == _T_643 ? $signed(7'sh10) : $signed(_GEN_18871); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18873 = 12'h6dd == _T_643 ? $signed(7'sh11) : $signed(_GEN_18872); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18874 = 12'h6de == _T_643 ? $signed(7'sh11) : $signed(_GEN_18873); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18875 = 12'h6df == _T_643 ? $signed(7'sh12) : $signed(_GEN_18874); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18876 = 12'h6e0 == _T_643 ? $signed(7'sh13) : $signed(_GEN_18875); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18877 = 12'h6e1 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18876); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18878 = 12'h6e2 == _T_643 ? $signed(7'sh14) : $signed(_GEN_18877); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18879 = 12'h6e3 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18878); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18880 = 12'h6e4 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18879); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18881 = 12'h6e5 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18880); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18882 = 12'h6e6 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18881); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18883 = 12'h6e7 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18882); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18884 = 12'h6e8 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18883); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18885 = 12'h6e9 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18884); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18886 = 12'h6ea == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18885); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18887 = 12'h6eb == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18886); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18888 = 12'h6ec == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18887); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18889 = 12'h6ed == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18888); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18890 = 12'h6ee == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18889); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18891 = 12'h6ef == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18890); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18892 = 12'h6f0 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18891); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18893 = 12'h6f1 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18892); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18894 = 12'h6f2 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18893); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18895 = 12'h6f3 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18894); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18896 = 12'h6f4 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18895); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18897 = 12'h6f5 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18896); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18898 = 12'h6f6 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18897); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18899 = 12'h6f7 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18898); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18900 = 12'h6f8 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18899); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18901 = 12'h6f9 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18900); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18902 = 12'h6fa == _T_643 ? $signed(7'sh25) : $signed(_GEN_18901); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18903 = 12'h6fb == _T_643 ? $signed(7'sh26) : $signed(_GEN_18902); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18904 = 12'h6fc == _T_643 ? $signed(7'sh27) : $signed(_GEN_18903); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18905 = 12'h6fd == _T_643 ? $signed(7'sh27) : $signed(_GEN_18904); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18906 = 12'h6fe == _T_643 ? $signed(7'sh28) : $signed(_GEN_18905); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18907 = 12'h6ff == _T_643 ? $signed(7'sh29) : $signed(_GEN_18906); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18908 = 12'h700 == _T_643 ? $signed(7'sh29) : $signed(_GEN_18907); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18909 = 12'h701 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_18908); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18910 = 12'h702 == _T_643 ? $signed(7'shb) : $signed(_GEN_18909); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18911 = 12'h703 == _T_643 ? $signed(7'shc) : $signed(_GEN_18910); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18912 = 12'h704 == _T_643 ? $signed(7'shc) : $signed(_GEN_18911); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18913 = 12'h705 == _T_643 ? $signed(7'shd) : $signed(_GEN_18912); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18914 = 12'h706 == _T_643 ? $signed(7'she) : $signed(_GEN_18913); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18915 = 12'h707 == _T_643 ? $signed(7'shf) : $signed(_GEN_18914); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18916 = 12'h708 == _T_643 ? $signed(7'shf) : $signed(_GEN_18915); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18917 = 12'h709 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18916); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18918 = 12'h70a == _T_643 ? $signed(7'sh11) : $signed(_GEN_18917); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18919 = 12'h70b == _T_643 ? $signed(7'sh11) : $signed(_GEN_18918); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18920 = 12'h70c == _T_643 ? $signed(7'sh12) : $signed(_GEN_18919); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18921 = 12'h70d == _T_643 ? $signed(7'sh13) : $signed(_GEN_18920); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18922 = 12'h70e == _T_643 ? $signed(7'sh14) : $signed(_GEN_18921); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18923 = 12'h70f == _T_643 ? $signed(7'sh14) : $signed(_GEN_18922); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18924 = 12'h710 == _T_643 ? $signed(7'sh15) : $signed(_GEN_18923); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18925 = 12'h711 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18924); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18926 = 12'h712 == _T_643 ? $signed(7'sh16) : $signed(_GEN_18925); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18927 = 12'h713 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18926); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18928 = 12'h714 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18927); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18929 = 12'h715 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18928); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18930 = 12'h716 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18929); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18931 = 12'h717 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18930); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18932 = 12'h718 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18931); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18933 = 12'h719 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18932); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18934 = 12'h71a == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18933); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18935 = 12'h71b == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18934); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18936 = 12'h71c == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18935); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18937 = 12'h71d == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18936); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18938 = 12'h71e == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18937); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18939 = 12'h71f == _T_643 ? $signed(7'sh20) : $signed(_GEN_18938); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18940 = 12'h720 == _T_643 ? $signed(7'sh20) : $signed(_GEN_18939); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18941 = 12'h721 == _T_643 ? $signed(7'sh21) : $signed(_GEN_18940); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18942 = 12'h722 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18941); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18943 = 12'h723 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18942); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18944 = 12'h724 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18943); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18945 = 12'h725 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18944); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18946 = 12'h726 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18945); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18947 = 12'h727 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18946); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18948 = 12'h728 == _T_643 ? $signed(7'sh26) : $signed(_GEN_18947); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18949 = 12'h729 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18948); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18950 = 12'h72a == _T_643 ? $signed(7'sh27) : $signed(_GEN_18949); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18951 = 12'h72b == _T_643 ? $signed(7'sh28) : $signed(_GEN_18950); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18952 = 12'h72c == _T_643 ? $signed(7'sh29) : $signed(_GEN_18951); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18953 = 12'h72d == _T_643 ? $signed(7'sh29) : $signed(_GEN_18952); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18954 = 12'h72e == _T_643 ? $signed(7'sh2a) : $signed(_GEN_18953); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18955 = 12'h72f == _T_643 ? $signed(7'sh2b) : $signed(_GEN_18954); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18956 = 12'h730 == _T_643 ? $signed(7'shc) : $signed(_GEN_18955); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18957 = 12'h731 == _T_643 ? $signed(7'shc) : $signed(_GEN_18956); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18958 = 12'h732 == _T_643 ? $signed(7'shd) : $signed(_GEN_18957); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18959 = 12'h733 == _T_643 ? $signed(7'she) : $signed(_GEN_18958); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18960 = 12'h734 == _T_643 ? $signed(7'shf) : $signed(_GEN_18959); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18961 = 12'h735 == _T_643 ? $signed(7'shf) : $signed(_GEN_18960); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18962 = 12'h736 == _T_643 ? $signed(7'sh10) : $signed(_GEN_18961); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18963 = 12'h737 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18962); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18964 = 12'h738 == _T_643 ? $signed(7'sh11) : $signed(_GEN_18963); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18965 = 12'h739 == _T_643 ? $signed(7'sh12) : $signed(_GEN_18964); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18966 = 12'h73a == _T_643 ? $signed(7'sh13) : $signed(_GEN_18965); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18967 = 12'h73b == _T_643 ? $signed(7'sh14) : $signed(_GEN_18966); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18968 = 12'h73c == _T_643 ? $signed(7'sh14) : $signed(_GEN_18967); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18969 = 12'h73d == _T_643 ? $signed(7'sh15) : $signed(_GEN_18968); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18970 = 12'h73e == _T_643 ? $signed(7'sh16) : $signed(_GEN_18969); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18971 = 12'h73f == _T_643 ? $signed(7'sh16) : $signed(_GEN_18970); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18972 = 12'h740 == _T_643 ? $signed(7'sh17) : $signed(_GEN_18971); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18973 = 12'h741 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18972); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18974 = 12'h742 == _T_643 ? $signed(7'sh18) : $signed(_GEN_18973); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18975 = 12'h743 == _T_643 ? $signed(7'sh19) : $signed(_GEN_18974); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18976 = 12'h744 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_18975); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18977 = 12'h745 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18976); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18978 = 12'h746 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_18977); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18979 = 12'h747 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_18978); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18980 = 12'h748 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18979); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18981 = 12'h749 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_18980); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18982 = 12'h74a == _T_643 ? $signed(7'sh1e) : $signed(_GEN_18981); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18983 = 12'h74b == _T_643 ? $signed(7'sh1f) : $signed(_GEN_18982); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18984 = 12'h74c == _T_643 ? $signed(7'sh20) : $signed(_GEN_18983); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18985 = 12'h74d == _T_643 ? $signed(7'sh20) : $signed(_GEN_18984); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18986 = 12'h74e == _T_643 ? $signed(7'sh21) : $signed(_GEN_18985); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18987 = 12'h74f == _T_643 ? $signed(7'sh22) : $signed(_GEN_18986); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18988 = 12'h750 == _T_643 ? $signed(7'sh22) : $signed(_GEN_18987); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18989 = 12'h751 == _T_643 ? $signed(7'sh23) : $signed(_GEN_18988); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18990 = 12'h752 == _T_643 ? $signed(7'sh24) : $signed(_GEN_18989); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18991 = 12'h753 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18990); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18992 = 12'h754 == _T_643 ? $signed(7'sh25) : $signed(_GEN_18991); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18993 = 12'h755 == _T_643 ? $signed(7'sh26) : $signed(_GEN_18992); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18994 = 12'h756 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18993); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18995 = 12'h757 == _T_643 ? $signed(7'sh27) : $signed(_GEN_18994); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18996 = 12'h758 == _T_643 ? $signed(7'sh28) : $signed(_GEN_18995); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18997 = 12'h759 == _T_643 ? $signed(7'sh29) : $signed(_GEN_18996); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18998 = 12'h75a == _T_643 ? $signed(7'sh29) : $signed(_GEN_18997); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_18999 = 12'h75b == _T_643 ? $signed(7'sh2a) : $signed(_GEN_18998); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19000 = 12'h75c == _T_643 ? $signed(7'sh2b) : $signed(_GEN_18999); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19001 = 12'h75d == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19000); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19002 = 12'h75e == _T_643 ? $signed(7'shc) : $signed(_GEN_19001); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19003 = 12'h75f == _T_643 ? $signed(7'shd) : $signed(_GEN_19002); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19004 = 12'h760 == _T_643 ? $signed(7'she) : $signed(_GEN_19003); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19005 = 12'h761 == _T_643 ? $signed(7'shf) : $signed(_GEN_19004); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19006 = 12'h762 == _T_643 ? $signed(7'shf) : $signed(_GEN_19005); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19007 = 12'h763 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19006); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19008 = 12'h764 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19007); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19009 = 12'h765 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19008); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19010 = 12'h766 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19009); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19011 = 12'h767 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19010); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19012 = 12'h768 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19011); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19013 = 12'h769 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19012); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19014 = 12'h76a == _T_643 ? $signed(7'sh15) : $signed(_GEN_19013); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19015 = 12'h76b == _T_643 ? $signed(7'sh16) : $signed(_GEN_19014); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19016 = 12'h76c == _T_643 ? $signed(7'sh16) : $signed(_GEN_19015); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19017 = 12'h76d == _T_643 ? $signed(7'sh17) : $signed(_GEN_19016); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19018 = 12'h76e == _T_643 ? $signed(7'sh18) : $signed(_GEN_19017); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19019 = 12'h76f == _T_643 ? $signed(7'sh18) : $signed(_GEN_19018); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19020 = 12'h770 == _T_643 ? $signed(7'sh19) : $signed(_GEN_19019); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19021 = 12'h771 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19020); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19022 = 12'h772 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19021); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19023 = 12'h773 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19022); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19024 = 12'h774 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_19023); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19025 = 12'h775 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19024); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19026 = 12'h776 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19025); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19027 = 12'h777 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_19026); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19028 = 12'h778 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_19027); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19029 = 12'h779 == _T_643 ? $signed(7'sh20) : $signed(_GEN_19028); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19030 = 12'h77a == _T_643 ? $signed(7'sh20) : $signed(_GEN_19029); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19031 = 12'h77b == _T_643 ? $signed(7'sh21) : $signed(_GEN_19030); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19032 = 12'h77c == _T_643 ? $signed(7'sh22) : $signed(_GEN_19031); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19033 = 12'h77d == _T_643 ? $signed(7'sh22) : $signed(_GEN_19032); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19034 = 12'h77e == _T_643 ? $signed(7'sh23) : $signed(_GEN_19033); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19035 = 12'h77f == _T_643 ? $signed(7'sh24) : $signed(_GEN_19034); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19036 = 12'h780 == _T_643 ? $signed(7'sh25) : $signed(_GEN_19035); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19037 = 12'h781 == _T_643 ? $signed(7'sh25) : $signed(_GEN_19036); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19038 = 12'h782 == _T_643 ? $signed(7'sh26) : $signed(_GEN_19037); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19039 = 12'h783 == _T_643 ? $signed(7'sh27) : $signed(_GEN_19038); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19040 = 12'h784 == _T_643 ? $signed(7'sh27) : $signed(_GEN_19039); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19041 = 12'h785 == _T_643 ? $signed(7'sh28) : $signed(_GEN_19040); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19042 = 12'h786 == _T_643 ? $signed(7'sh29) : $signed(_GEN_19041); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19043 = 12'h787 == _T_643 ? $signed(7'sh29) : $signed(_GEN_19042); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19044 = 12'h788 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_19043); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19045 = 12'h789 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_19044); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19046 = 12'h78a == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19045); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19047 = 12'h78b == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19046); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19048 = 12'h78c == _T_643 ? $signed(7'shd) : $signed(_GEN_19047); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19049 = 12'h78d == _T_643 ? $signed(7'she) : $signed(_GEN_19048); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19050 = 12'h78e == _T_643 ? $signed(7'shf) : $signed(_GEN_19049); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19051 = 12'h78f == _T_643 ? $signed(7'shf) : $signed(_GEN_19050); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19052 = 12'h790 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19051); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19053 = 12'h791 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19052); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19054 = 12'h792 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19053); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19055 = 12'h793 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19054); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19056 = 12'h794 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19055); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19057 = 12'h795 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19056); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19058 = 12'h796 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19057); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19059 = 12'h797 == _T_643 ? $signed(7'sh15) : $signed(_GEN_19058); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19060 = 12'h798 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19059); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19061 = 12'h799 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19060); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19062 = 12'h79a == _T_643 ? $signed(7'sh17) : $signed(_GEN_19061); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19063 = 12'h79b == _T_643 ? $signed(7'sh18) : $signed(_GEN_19062); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19064 = 12'h79c == _T_643 ? $signed(7'sh18) : $signed(_GEN_19063); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19065 = 12'h79d == _T_643 ? $signed(7'sh19) : $signed(_GEN_19064); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19066 = 12'h79e == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19065); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19067 = 12'h79f == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19066); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19068 = 12'h7a0 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19067); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19069 = 12'h7a1 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_19068); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19070 = 12'h7a2 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19069); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19071 = 12'h7a3 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19070); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19072 = 12'h7a4 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_19071); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19073 = 12'h7a5 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_19072); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19074 = 12'h7a6 == _T_643 ? $signed(7'sh20) : $signed(_GEN_19073); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19075 = 12'h7a7 == _T_643 ? $signed(7'sh20) : $signed(_GEN_19074); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19076 = 12'h7a8 == _T_643 ? $signed(7'sh21) : $signed(_GEN_19075); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19077 = 12'h7a9 == _T_643 ? $signed(7'sh22) : $signed(_GEN_19076); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19078 = 12'h7aa == _T_643 ? $signed(7'sh22) : $signed(_GEN_19077); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19079 = 12'h7ab == _T_643 ? $signed(7'sh23) : $signed(_GEN_19078); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19080 = 12'h7ac == _T_643 ? $signed(7'sh24) : $signed(_GEN_19079); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19081 = 12'h7ad == _T_643 ? $signed(7'sh25) : $signed(_GEN_19080); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19082 = 12'h7ae == _T_643 ? $signed(7'sh25) : $signed(_GEN_19081); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19083 = 12'h7af == _T_643 ? $signed(7'sh26) : $signed(_GEN_19082); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19084 = 12'h7b0 == _T_643 ? $signed(7'sh27) : $signed(_GEN_19083); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19085 = 12'h7b1 == _T_643 ? $signed(7'sh27) : $signed(_GEN_19084); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19086 = 12'h7b2 == _T_643 ? $signed(7'sh28) : $signed(_GEN_19085); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19087 = 12'h7b3 == _T_643 ? $signed(7'sh29) : $signed(_GEN_19086); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19088 = 12'h7b4 == _T_643 ? $signed(7'sh29) : $signed(_GEN_19087); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19089 = 12'h7b5 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_19088); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19090 = 12'h7b6 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_19089); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19091 = 12'h7b7 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19090); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19092 = 12'h7b8 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19091); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19093 = 12'h7b9 == _T_643 ? $signed(7'sh2d) : $signed(_GEN_19092); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19094 = 12'h7ba == _T_643 ? $signed(7'she) : $signed(_GEN_19093); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19095 = 12'h7bb == _T_643 ? $signed(7'shf) : $signed(_GEN_19094); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19096 = 12'h7bc == _T_643 ? $signed(7'shf) : $signed(_GEN_19095); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19097 = 12'h7bd == _T_643 ? $signed(7'sh10) : $signed(_GEN_19096); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19098 = 12'h7be == _T_643 ? $signed(7'sh11) : $signed(_GEN_19097); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19099 = 12'h7bf == _T_643 ? $signed(7'sh11) : $signed(_GEN_19098); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19100 = 12'h7c0 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19099); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19101 = 12'h7c1 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19100); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19102 = 12'h7c2 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19101); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19103 = 12'h7c3 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19102); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19104 = 12'h7c4 == _T_643 ? $signed(7'sh15) : $signed(_GEN_19103); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19105 = 12'h7c5 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19104); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19106 = 12'h7c6 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19105); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19107 = 12'h7c7 == _T_643 ? $signed(7'sh17) : $signed(_GEN_19106); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19108 = 12'h7c8 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19107); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19109 = 12'h7c9 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19108); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19110 = 12'h7ca == _T_643 ? $signed(7'sh19) : $signed(_GEN_19109); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19111 = 12'h7cb == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19110); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19112 = 12'h7cc == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19111); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19113 = 12'h7cd == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19112); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19114 = 12'h7ce == _T_643 ? $signed(7'sh1c) : $signed(_GEN_19113); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19115 = 12'h7cf == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19114); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19116 = 12'h7d0 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19115); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19117 = 12'h7d1 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_19116); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19118 = 12'h7d2 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_19117); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19119 = 12'h7d3 == _T_643 ? $signed(7'sh20) : $signed(_GEN_19118); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19120 = 12'h7d4 == _T_643 ? $signed(7'sh20) : $signed(_GEN_19119); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19121 = 12'h7d5 == _T_643 ? $signed(7'sh21) : $signed(_GEN_19120); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19122 = 12'h7d6 == _T_643 ? $signed(7'sh22) : $signed(_GEN_19121); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19123 = 12'h7d7 == _T_643 ? $signed(7'sh22) : $signed(_GEN_19122); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19124 = 12'h7d8 == _T_643 ? $signed(7'sh23) : $signed(_GEN_19123); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19125 = 12'h7d9 == _T_643 ? $signed(7'sh24) : $signed(_GEN_19124); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19126 = 12'h7da == _T_643 ? $signed(7'sh25) : $signed(_GEN_19125); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19127 = 12'h7db == _T_643 ? $signed(7'sh25) : $signed(_GEN_19126); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19128 = 12'h7dc == _T_643 ? $signed(7'sh26) : $signed(_GEN_19127); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19129 = 12'h7dd == _T_643 ? $signed(7'sh27) : $signed(_GEN_19128); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19130 = 12'h7de == _T_643 ? $signed(7'sh27) : $signed(_GEN_19129); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19131 = 12'h7df == _T_643 ? $signed(7'sh28) : $signed(_GEN_19130); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19132 = 12'h7e0 == _T_643 ? $signed(7'sh29) : $signed(_GEN_19131); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19133 = 12'h7e1 == _T_643 ? $signed(7'sh29) : $signed(_GEN_19132); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19134 = 12'h7e2 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_19133); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19135 = 12'h7e3 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_19134); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19136 = 12'h7e4 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19135); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19137 = 12'h7e5 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19136); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19138 = 12'h7e6 == _T_643 ? $signed(7'sh2d) : $signed(_GEN_19137); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19139 = 12'h7e7 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_19138); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19140 = 12'h7e8 == _T_643 ? $signed(7'shf) : $signed(_GEN_19139); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19141 = 12'h7e9 == _T_643 ? $signed(7'shf) : $signed(_GEN_19140); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19142 = 12'h7ea == _T_643 ? $signed(7'sh10) : $signed(_GEN_19141); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19143 = 12'h7eb == _T_643 ? $signed(7'sh11) : $signed(_GEN_19142); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19144 = 12'h7ec == _T_643 ? $signed(7'sh11) : $signed(_GEN_19143); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19145 = 12'h7ed == _T_643 ? $signed(7'sh12) : $signed(_GEN_19144); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19146 = 12'h7ee == _T_643 ? $signed(7'sh13) : $signed(_GEN_19145); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19147 = 12'h7ef == _T_643 ? $signed(7'sh14) : $signed(_GEN_19146); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19148 = 12'h7f0 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19147); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19149 = 12'h7f1 == _T_643 ? $signed(7'sh15) : $signed(_GEN_19148); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19150 = 12'h7f2 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19149); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19151 = 12'h7f3 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19150); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19152 = 12'h7f4 == _T_643 ? $signed(7'sh17) : $signed(_GEN_19151); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19153 = 12'h7f5 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19152); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19154 = 12'h7f6 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19153); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19155 = 12'h7f7 == _T_643 ? $signed(7'sh19) : $signed(_GEN_19154); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19156 = 12'h7f8 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19155); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19157 = 12'h7f9 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19156); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19158 = 12'h7fa == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19157); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19159 = 12'h7fb == _T_643 ? $signed(7'sh1c) : $signed(_GEN_19158); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19160 = 12'h7fc == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19159); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19161 = 12'h7fd == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19160); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19162 = 12'h7fe == _T_643 ? $signed(7'sh1e) : $signed(_GEN_19161); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19163 = 12'h7ff == _T_643 ? $signed(7'sh1f) : $signed(_GEN_19162); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19164 = 12'h800 == _T_643 ? $signed(7'sh20) : $signed(_GEN_19163); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19165 = 12'h801 == _T_643 ? $signed(7'sh20) : $signed(_GEN_19164); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19166 = 12'h802 == _T_643 ? $signed(7'sh21) : $signed(_GEN_19165); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19167 = 12'h803 == _T_643 ? $signed(7'sh22) : $signed(_GEN_19166); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19168 = 12'h804 == _T_643 ? $signed(7'sh22) : $signed(_GEN_19167); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19169 = 12'h805 == _T_643 ? $signed(7'sh23) : $signed(_GEN_19168); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19170 = 12'h806 == _T_643 ? $signed(7'sh24) : $signed(_GEN_19169); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19171 = 12'h807 == _T_643 ? $signed(7'sh25) : $signed(_GEN_19170); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19172 = 12'h808 == _T_643 ? $signed(7'sh25) : $signed(_GEN_19171); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19173 = 12'h809 == _T_643 ? $signed(7'sh26) : $signed(_GEN_19172); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19174 = 12'h80a == _T_643 ? $signed(7'sh27) : $signed(_GEN_19173); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19175 = 12'h80b == _T_643 ? $signed(7'sh27) : $signed(_GEN_19174); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19176 = 12'h80c == _T_643 ? $signed(7'sh28) : $signed(_GEN_19175); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19177 = 12'h80d == _T_643 ? $signed(7'sh29) : $signed(_GEN_19176); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19178 = 12'h80e == _T_643 ? $signed(7'sh29) : $signed(_GEN_19177); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19179 = 12'h80f == _T_643 ? $signed(7'sh2a) : $signed(_GEN_19178); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19180 = 12'h810 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_19179); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19181 = 12'h811 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19180); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19182 = 12'h812 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19181); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19183 = 12'h813 == _T_643 ? $signed(7'sh2d) : $signed(_GEN_19182); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19184 = 12'h814 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_19183); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19185 = 12'h815 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_19184); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19186 = 12'h816 == _T_643 ? $signed(7'shf) : $signed(_GEN_19185); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19187 = 12'h817 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19186); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19188 = 12'h818 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19187); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19189 = 12'h819 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19188); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19190 = 12'h81a == _T_643 ? $signed(7'sh12) : $signed(_GEN_19189); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19191 = 12'h81b == _T_643 ? $signed(7'sh13) : $signed(_GEN_19190); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19192 = 12'h81c == _T_643 ? $signed(7'sh14) : $signed(_GEN_19191); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19193 = 12'h81d == _T_643 ? $signed(7'sh14) : $signed(_GEN_19192); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19194 = 12'h81e == _T_643 ? $signed(7'sh15) : $signed(_GEN_19193); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19195 = 12'h81f == _T_643 ? $signed(7'sh16) : $signed(_GEN_19194); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19196 = 12'h820 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19195); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19197 = 12'h821 == _T_643 ? $signed(7'sh17) : $signed(_GEN_19196); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19198 = 12'h822 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19197); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19199 = 12'h823 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19198); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19200 = 12'h824 == _T_643 ? $signed(7'sh19) : $signed(_GEN_19199); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19201 = 12'h825 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19200); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19202 = 12'h826 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19201); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19203 = 12'h827 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19202); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19204 = 12'h828 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_19203); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19205 = 12'h829 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19204); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19206 = 12'h82a == _T_643 ? $signed(7'sh1d) : $signed(_GEN_19205); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19207 = 12'h82b == _T_643 ? $signed(7'sh1e) : $signed(_GEN_19206); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19208 = 12'h82c == _T_643 ? $signed(7'sh1f) : $signed(_GEN_19207); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19209 = 12'h82d == _T_643 ? $signed(7'sh20) : $signed(_GEN_19208); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19210 = 12'h82e == _T_643 ? $signed(7'sh20) : $signed(_GEN_19209); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19211 = 12'h82f == _T_643 ? $signed(7'sh21) : $signed(_GEN_19210); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19212 = 12'h830 == _T_643 ? $signed(7'sh22) : $signed(_GEN_19211); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19213 = 12'h831 == _T_643 ? $signed(7'sh22) : $signed(_GEN_19212); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19214 = 12'h832 == _T_643 ? $signed(7'sh23) : $signed(_GEN_19213); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19215 = 12'h833 == _T_643 ? $signed(7'sh24) : $signed(_GEN_19214); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19216 = 12'h834 == _T_643 ? $signed(7'sh25) : $signed(_GEN_19215); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19217 = 12'h835 == _T_643 ? $signed(7'sh25) : $signed(_GEN_19216); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19218 = 12'h836 == _T_643 ? $signed(7'sh26) : $signed(_GEN_19217); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19219 = 12'h837 == _T_643 ? $signed(7'sh27) : $signed(_GEN_19218); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19220 = 12'h838 == _T_643 ? $signed(7'sh27) : $signed(_GEN_19219); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19221 = 12'h839 == _T_643 ? $signed(7'sh28) : $signed(_GEN_19220); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19222 = 12'h83a == _T_643 ? $signed(7'sh29) : $signed(_GEN_19221); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19223 = 12'h83b == _T_643 ? $signed(7'sh29) : $signed(_GEN_19222); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19224 = 12'h83c == _T_643 ? $signed(7'sh2a) : $signed(_GEN_19223); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19225 = 12'h83d == _T_643 ? $signed(7'sh2b) : $signed(_GEN_19224); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19226 = 12'h83e == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19225); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19227 = 12'h83f == _T_643 ? $signed(7'sh2c) : $signed(_GEN_19226); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19228 = 12'h840 == _T_643 ? $signed(7'sh2d) : $signed(_GEN_19227); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19229 = 12'h841 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_19228); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19230 = 12'h842 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_19229); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19231 = 12'h843 == _T_643 ? $signed(7'sh2f) : $signed(_GEN_19230); // @[GraphicEngineVGA.scala 321:24]
  wire [11:0] inSpriteX_4 = spriteRotationReg_4 ? $signed({{5{_GEN_19231[6]}},_GEN_19231}) : $signed(_T_628); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_19233 = 12'h1 == _T_643 ? $signed(7'shf) : $signed(7'sh10); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19234 = 12'h2 == _T_643 ? $signed(7'shf) : $signed(_GEN_19233); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19235 = 12'h3 == _T_643 ? $signed(7'she) : $signed(_GEN_19234); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19236 = 12'h4 == _T_643 ? $signed(7'shd) : $signed(_GEN_19235); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19237 = 12'h5 == _T_643 ? $signed(7'shc) : $signed(_GEN_19236); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19238 = 12'h6 == _T_643 ? $signed(7'shc) : $signed(_GEN_19237); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19239 = 12'h7 == _T_643 ? $signed(7'shb) : $signed(_GEN_19238); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19240 = 12'h8 == _T_643 ? $signed(7'sha) : $signed(_GEN_19239); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19241 = 12'h9 == _T_643 ? $signed(7'sha) : $signed(_GEN_19240); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19242 = 12'ha == _T_643 ? $signed(7'sh9) : $signed(_GEN_19241); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19243 = 12'hb == _T_643 ? $signed(7'sh8) : $signed(_GEN_19242); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19244 = 12'hc == _T_643 ? $signed(7'sh8) : $signed(_GEN_19243); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19245 = 12'hd == _T_643 ? $signed(7'sh7) : $signed(_GEN_19244); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19246 = 12'he == _T_643 ? $signed(7'sh6) : $signed(_GEN_19245); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19247 = 12'hf == _T_643 ? $signed(7'sh5) : $signed(_GEN_19246); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19248 = 12'h10 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19247); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19249 = 12'h11 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19248); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19250 = 12'h12 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19249); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19251 = 12'h13 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19250); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19252 = 12'h14 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19251); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19253 = 12'h15 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19252); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19254 = 12'h16 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19253); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19255 = 12'h17 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19254); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19256 = 12'h18 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19255); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19257 = 12'h19 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19256); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19258 = 12'h1a == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19257); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19259 = 12'h1b == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19258); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19260 = 12'h1c == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19259); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19261 = 12'h1d == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19260); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19262 = 12'h1e == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19261); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19263 = 12'h1f == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19262); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19264 = 12'h20 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19263); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19265 = 12'h21 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19264); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19266 = 12'h22 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19265); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19267 = 12'h23 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19266); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19268 = 12'h24 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19267); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19269 = 12'h25 == _T_643 ? $signed(-7'sha) : $signed(_GEN_19268); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19270 = 12'h26 == _T_643 ? $signed(-7'shb) : $signed(_GEN_19269); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19271 = 12'h27 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19270); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19272 = 12'h28 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19271); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19273 = 12'h29 == _T_643 ? $signed(-7'shd) : $signed(_GEN_19272); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19274 = 12'h2a == _T_643 ? $signed(-7'she) : $signed(_GEN_19273); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19275 = 12'h2b == _T_643 ? $signed(-7'she) : $signed(_GEN_19274); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19276 = 12'h2c == _T_643 ? $signed(-7'shf) : $signed(_GEN_19275); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19277 = 12'h2d == _T_643 ? $signed(-7'sh10) : $signed(_GEN_19276); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19278 = 12'h2e == _T_643 ? $signed(7'sh11) : $signed(_GEN_19277); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19279 = 12'h2f == _T_643 ? $signed(7'sh10) : $signed(_GEN_19278); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19280 = 12'h30 == _T_643 ? $signed(7'shf) : $signed(_GEN_19279); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19281 = 12'h31 == _T_643 ? $signed(7'shf) : $signed(_GEN_19280); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19282 = 12'h32 == _T_643 ? $signed(7'she) : $signed(_GEN_19281); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19283 = 12'h33 == _T_643 ? $signed(7'shd) : $signed(_GEN_19282); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19284 = 12'h34 == _T_643 ? $signed(7'shc) : $signed(_GEN_19283); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19285 = 12'h35 == _T_643 ? $signed(7'shc) : $signed(_GEN_19284); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19286 = 12'h36 == _T_643 ? $signed(7'shb) : $signed(_GEN_19285); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19287 = 12'h37 == _T_643 ? $signed(7'sha) : $signed(_GEN_19286); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19288 = 12'h38 == _T_643 ? $signed(7'sha) : $signed(_GEN_19287); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19289 = 12'h39 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19288); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19290 = 12'h3a == _T_643 ? $signed(7'sh8) : $signed(_GEN_19289); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19291 = 12'h3b == _T_643 ? $signed(7'sh8) : $signed(_GEN_19290); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19292 = 12'h3c == _T_643 ? $signed(7'sh7) : $signed(_GEN_19291); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19293 = 12'h3d == _T_643 ? $signed(7'sh6) : $signed(_GEN_19292); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19294 = 12'h3e == _T_643 ? $signed(7'sh5) : $signed(_GEN_19293); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19295 = 12'h3f == _T_643 ? $signed(7'sh5) : $signed(_GEN_19294); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19296 = 12'h40 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19295); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19297 = 12'h41 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19296); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19298 = 12'h42 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19297); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19299 = 12'h43 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19298); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19300 = 12'h44 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19299); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19301 = 12'h45 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19300); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19302 = 12'h46 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19301); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19303 = 12'h47 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19302); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19304 = 12'h48 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19303); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19305 = 12'h49 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19304); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19306 = 12'h4a == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19305); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19307 = 12'h4b == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19306); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19308 = 12'h4c == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19307); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19309 = 12'h4d == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19308); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19310 = 12'h4e == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19309); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19311 = 12'h4f == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19310); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19312 = 12'h50 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19311); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19313 = 12'h51 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19312); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19314 = 12'h52 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19313); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19315 = 12'h53 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19314); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19316 = 12'h54 == _T_643 ? $signed(-7'sha) : $signed(_GEN_19315); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19317 = 12'h55 == _T_643 ? $signed(-7'shb) : $signed(_GEN_19316); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19318 = 12'h56 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19317); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19319 = 12'h57 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19318); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19320 = 12'h58 == _T_643 ? $signed(-7'shd) : $signed(_GEN_19319); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19321 = 12'h59 == _T_643 ? $signed(-7'she) : $signed(_GEN_19320); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19322 = 12'h5a == _T_643 ? $signed(-7'she) : $signed(_GEN_19321); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19323 = 12'h5b == _T_643 ? $signed(-7'shf) : $signed(_GEN_19322); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19324 = 12'h5c == _T_643 ? $signed(7'sh11) : $signed(_GEN_19323); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19325 = 12'h5d == _T_643 ? $signed(7'sh11) : $signed(_GEN_19324); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19326 = 12'h5e == _T_643 ? $signed(7'sh10) : $signed(_GEN_19325); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19327 = 12'h5f == _T_643 ? $signed(7'shf) : $signed(_GEN_19326); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19328 = 12'h60 == _T_643 ? $signed(7'shf) : $signed(_GEN_19327); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19329 = 12'h61 == _T_643 ? $signed(7'she) : $signed(_GEN_19328); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19330 = 12'h62 == _T_643 ? $signed(7'shd) : $signed(_GEN_19329); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19331 = 12'h63 == _T_643 ? $signed(7'shc) : $signed(_GEN_19330); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19332 = 12'h64 == _T_643 ? $signed(7'shc) : $signed(_GEN_19331); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19333 = 12'h65 == _T_643 ? $signed(7'shb) : $signed(_GEN_19332); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19334 = 12'h66 == _T_643 ? $signed(7'sha) : $signed(_GEN_19333); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19335 = 12'h67 == _T_643 ? $signed(7'sha) : $signed(_GEN_19334); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19336 = 12'h68 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19335); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19337 = 12'h69 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19336); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19338 = 12'h6a == _T_643 ? $signed(7'sh8) : $signed(_GEN_19337); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19339 = 12'h6b == _T_643 ? $signed(7'sh7) : $signed(_GEN_19338); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19340 = 12'h6c == _T_643 ? $signed(7'sh6) : $signed(_GEN_19339); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19341 = 12'h6d == _T_643 ? $signed(7'sh5) : $signed(_GEN_19340); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19342 = 12'h6e == _T_643 ? $signed(7'sh5) : $signed(_GEN_19341); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19343 = 12'h6f == _T_643 ? $signed(7'sh4) : $signed(_GEN_19342); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19344 = 12'h70 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19343); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19345 = 12'h71 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19344); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19346 = 12'h72 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19345); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19347 = 12'h73 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19346); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19348 = 12'h74 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19347); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19349 = 12'h75 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19348); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19350 = 12'h76 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19349); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19351 = 12'h77 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19350); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19352 = 12'h78 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19351); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19353 = 12'h79 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19352); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19354 = 12'h7a == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19353); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19355 = 12'h7b == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19354); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19356 = 12'h7c == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19355); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19357 = 12'h7d == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19356); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19358 = 12'h7e == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19357); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19359 = 12'h7f == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19358); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19360 = 12'h80 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19359); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19361 = 12'h81 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19360); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19362 = 12'h82 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19361); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19363 = 12'h83 == _T_643 ? $signed(-7'sha) : $signed(_GEN_19362); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19364 = 12'h84 == _T_643 ? $signed(-7'shb) : $signed(_GEN_19363); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19365 = 12'h85 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19364); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19366 = 12'h86 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19365); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19367 = 12'h87 == _T_643 ? $signed(-7'shd) : $signed(_GEN_19366); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19368 = 12'h88 == _T_643 ? $signed(-7'she) : $signed(_GEN_19367); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19369 = 12'h89 == _T_643 ? $signed(-7'she) : $signed(_GEN_19368); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19370 = 12'h8a == _T_643 ? $signed(7'sh12) : $signed(_GEN_19369); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19371 = 12'h8b == _T_643 ? $signed(7'sh11) : $signed(_GEN_19370); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19372 = 12'h8c == _T_643 ? $signed(7'sh11) : $signed(_GEN_19371); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19373 = 12'h8d == _T_643 ? $signed(7'sh10) : $signed(_GEN_19372); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19374 = 12'h8e == _T_643 ? $signed(7'shf) : $signed(_GEN_19373); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19375 = 12'h8f == _T_643 ? $signed(7'shf) : $signed(_GEN_19374); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19376 = 12'h90 == _T_643 ? $signed(7'she) : $signed(_GEN_19375); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19377 = 12'h91 == _T_643 ? $signed(7'shd) : $signed(_GEN_19376); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19378 = 12'h92 == _T_643 ? $signed(7'shc) : $signed(_GEN_19377); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19379 = 12'h93 == _T_643 ? $signed(7'shc) : $signed(_GEN_19378); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19380 = 12'h94 == _T_643 ? $signed(7'shb) : $signed(_GEN_19379); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19381 = 12'h95 == _T_643 ? $signed(7'sha) : $signed(_GEN_19380); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19382 = 12'h96 == _T_643 ? $signed(7'sha) : $signed(_GEN_19381); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19383 = 12'h97 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19382); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19384 = 12'h98 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19383); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19385 = 12'h99 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19384); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19386 = 12'h9a == _T_643 ? $signed(7'sh7) : $signed(_GEN_19385); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19387 = 12'h9b == _T_643 ? $signed(7'sh6) : $signed(_GEN_19386); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19388 = 12'h9c == _T_643 ? $signed(7'sh5) : $signed(_GEN_19387); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19389 = 12'h9d == _T_643 ? $signed(7'sh5) : $signed(_GEN_19388); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19390 = 12'h9e == _T_643 ? $signed(7'sh4) : $signed(_GEN_19389); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19391 = 12'h9f == _T_643 ? $signed(7'sh3) : $signed(_GEN_19390); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19392 = 12'ha0 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19391); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19393 = 12'ha1 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19392); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19394 = 12'ha2 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19393); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19395 = 12'ha3 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19394); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19396 = 12'ha4 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19395); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19397 = 12'ha5 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19396); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19398 = 12'ha6 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19397); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19399 = 12'ha7 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19398); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19400 = 12'ha8 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19399); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19401 = 12'ha9 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19400); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19402 = 12'haa == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19401); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19403 = 12'hab == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19402); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19404 = 12'hac == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19403); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19405 = 12'had == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19404); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19406 = 12'hae == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19405); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19407 = 12'haf == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19406); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19408 = 12'hb0 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19407); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19409 = 12'hb1 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19408); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19410 = 12'hb2 == _T_643 ? $signed(-7'sha) : $signed(_GEN_19409); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19411 = 12'hb3 == _T_643 ? $signed(-7'shb) : $signed(_GEN_19410); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19412 = 12'hb4 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19411); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19413 = 12'hb5 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19412); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19414 = 12'hb6 == _T_643 ? $signed(-7'shd) : $signed(_GEN_19413); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19415 = 12'hb7 == _T_643 ? $signed(-7'she) : $signed(_GEN_19414); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19416 = 12'hb8 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19415); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19417 = 12'hb9 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19416); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19418 = 12'hba == _T_643 ? $signed(7'sh11) : $signed(_GEN_19417); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19419 = 12'hbb == _T_643 ? $signed(7'sh11) : $signed(_GEN_19418); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19420 = 12'hbc == _T_643 ? $signed(7'sh10) : $signed(_GEN_19419); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19421 = 12'hbd == _T_643 ? $signed(7'shf) : $signed(_GEN_19420); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19422 = 12'hbe == _T_643 ? $signed(7'shf) : $signed(_GEN_19421); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19423 = 12'hbf == _T_643 ? $signed(7'she) : $signed(_GEN_19422); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19424 = 12'hc0 == _T_643 ? $signed(7'shd) : $signed(_GEN_19423); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19425 = 12'hc1 == _T_643 ? $signed(7'shc) : $signed(_GEN_19424); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19426 = 12'hc2 == _T_643 ? $signed(7'shc) : $signed(_GEN_19425); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19427 = 12'hc3 == _T_643 ? $signed(7'shb) : $signed(_GEN_19426); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19428 = 12'hc4 == _T_643 ? $signed(7'sha) : $signed(_GEN_19427); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19429 = 12'hc5 == _T_643 ? $signed(7'sha) : $signed(_GEN_19428); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19430 = 12'hc6 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19429); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19431 = 12'hc7 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19430); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19432 = 12'hc8 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19431); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19433 = 12'hc9 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19432); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19434 = 12'hca == _T_643 ? $signed(7'sh6) : $signed(_GEN_19433); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19435 = 12'hcb == _T_643 ? $signed(7'sh5) : $signed(_GEN_19434); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19436 = 12'hcc == _T_643 ? $signed(7'sh5) : $signed(_GEN_19435); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19437 = 12'hcd == _T_643 ? $signed(7'sh4) : $signed(_GEN_19436); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19438 = 12'hce == _T_643 ? $signed(7'sh3) : $signed(_GEN_19437); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19439 = 12'hcf == _T_643 ? $signed(7'sh3) : $signed(_GEN_19438); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19440 = 12'hd0 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19439); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19441 = 12'hd1 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19440); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19442 = 12'hd2 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19441); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19443 = 12'hd3 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19442); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19444 = 12'hd4 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19443); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19445 = 12'hd5 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19444); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19446 = 12'hd6 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19445); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19447 = 12'hd7 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19446); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19448 = 12'hd8 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19447); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19449 = 12'hd9 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19448); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19450 = 12'hda == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19449); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19451 = 12'hdb == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19450); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19452 = 12'hdc == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19451); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19453 = 12'hdd == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19452); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19454 = 12'hde == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19453); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19455 = 12'hdf == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19454); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19456 = 12'he0 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19455); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19457 = 12'he1 == _T_643 ? $signed(-7'sha) : $signed(_GEN_19456); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19458 = 12'he2 == _T_643 ? $signed(-7'shb) : $signed(_GEN_19457); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19459 = 12'he3 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19458); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19460 = 12'he4 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19459); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19461 = 12'he5 == _T_643 ? $signed(-7'shd) : $signed(_GEN_19460); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19462 = 12'he6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19461); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19463 = 12'he7 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19462); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19464 = 12'he8 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19463); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19465 = 12'he9 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19464); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19466 = 12'hea == _T_643 ? $signed(7'sh11) : $signed(_GEN_19465); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19467 = 12'heb == _T_643 ? $signed(7'sh10) : $signed(_GEN_19466); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19468 = 12'hec == _T_643 ? $signed(7'shf) : $signed(_GEN_19467); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19469 = 12'hed == _T_643 ? $signed(7'shf) : $signed(_GEN_19468); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19470 = 12'hee == _T_643 ? $signed(7'she) : $signed(_GEN_19469); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19471 = 12'hef == _T_643 ? $signed(7'shd) : $signed(_GEN_19470); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19472 = 12'hf0 == _T_643 ? $signed(7'shc) : $signed(_GEN_19471); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19473 = 12'hf1 == _T_643 ? $signed(7'shc) : $signed(_GEN_19472); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19474 = 12'hf2 == _T_643 ? $signed(7'shb) : $signed(_GEN_19473); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19475 = 12'hf3 == _T_643 ? $signed(7'sha) : $signed(_GEN_19474); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19476 = 12'hf4 == _T_643 ? $signed(7'sha) : $signed(_GEN_19475); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19477 = 12'hf5 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19476); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19478 = 12'hf6 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19477); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19479 = 12'hf7 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19478); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19480 = 12'hf8 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19479); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19481 = 12'hf9 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19480); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19482 = 12'hfa == _T_643 ? $signed(7'sh5) : $signed(_GEN_19481); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19483 = 12'hfb == _T_643 ? $signed(7'sh5) : $signed(_GEN_19482); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19484 = 12'hfc == _T_643 ? $signed(7'sh4) : $signed(_GEN_19483); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19485 = 12'hfd == _T_643 ? $signed(7'sh3) : $signed(_GEN_19484); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19486 = 12'hfe == _T_643 ? $signed(7'sh3) : $signed(_GEN_19485); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19487 = 12'hff == _T_643 ? $signed(7'sh2) : $signed(_GEN_19486); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19488 = 12'h100 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19487); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19489 = 12'h101 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19488); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19490 = 12'h102 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19489); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19491 = 12'h103 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19490); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19492 = 12'h104 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19491); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19493 = 12'h105 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19492); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19494 = 12'h106 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19493); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19495 = 12'h107 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19494); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19496 = 12'h108 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19495); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19497 = 12'h109 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19496); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19498 = 12'h10a == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19497); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19499 = 12'h10b == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19498); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19500 = 12'h10c == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19499); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19501 = 12'h10d == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19500); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19502 = 12'h10e == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19501); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19503 = 12'h10f == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19502); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19504 = 12'h110 == _T_643 ? $signed(-7'sha) : $signed(_GEN_19503); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19505 = 12'h111 == _T_643 ? $signed(-7'shb) : $signed(_GEN_19504); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19506 = 12'h112 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19505); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19507 = 12'h113 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19506); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19508 = 12'h114 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19507); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19509 = 12'h115 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19508); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19510 = 12'h116 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19509); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19511 = 12'h117 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19510); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19512 = 12'h118 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19511); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19513 = 12'h119 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19512); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19514 = 12'h11a == _T_643 ? $signed(7'sh10) : $signed(_GEN_19513); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19515 = 12'h11b == _T_643 ? $signed(7'shf) : $signed(_GEN_19514); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19516 = 12'h11c == _T_643 ? $signed(7'shf) : $signed(_GEN_19515); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19517 = 12'h11d == _T_643 ? $signed(7'she) : $signed(_GEN_19516); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19518 = 12'h11e == _T_643 ? $signed(7'shd) : $signed(_GEN_19517); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19519 = 12'h11f == _T_643 ? $signed(7'shc) : $signed(_GEN_19518); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19520 = 12'h120 == _T_643 ? $signed(7'shc) : $signed(_GEN_19519); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19521 = 12'h121 == _T_643 ? $signed(7'shb) : $signed(_GEN_19520); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19522 = 12'h122 == _T_643 ? $signed(7'sha) : $signed(_GEN_19521); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19523 = 12'h123 == _T_643 ? $signed(7'sha) : $signed(_GEN_19522); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19524 = 12'h124 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19523); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19525 = 12'h125 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19524); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19526 = 12'h126 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19525); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19527 = 12'h127 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19526); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19528 = 12'h128 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19527); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19529 = 12'h129 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19528); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19530 = 12'h12a == _T_643 ? $signed(7'sh5) : $signed(_GEN_19529); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19531 = 12'h12b == _T_643 ? $signed(7'sh4) : $signed(_GEN_19530); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19532 = 12'h12c == _T_643 ? $signed(7'sh3) : $signed(_GEN_19531); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19533 = 12'h12d == _T_643 ? $signed(7'sh3) : $signed(_GEN_19532); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19534 = 12'h12e == _T_643 ? $signed(7'sh2) : $signed(_GEN_19533); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19535 = 12'h12f == _T_643 ? $signed(7'sh1) : $signed(_GEN_19534); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19536 = 12'h130 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19535); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19537 = 12'h131 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19536); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19538 = 12'h132 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19537); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19539 = 12'h133 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19538); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19540 = 12'h134 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19539); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19541 = 12'h135 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19540); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19542 = 12'h136 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19541); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19543 = 12'h137 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19542); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19544 = 12'h138 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19543); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19545 = 12'h139 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19544); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19546 = 12'h13a == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19545); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19547 = 12'h13b == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19546); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19548 = 12'h13c == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19547); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19549 = 12'h13d == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19548); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19550 = 12'h13e == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19549); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19551 = 12'h13f == _T_643 ? $signed(-7'sha) : $signed(_GEN_19550); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19552 = 12'h140 == _T_643 ? $signed(-7'shb) : $signed(_GEN_19551); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19553 = 12'h141 == _T_643 ? $signed(-7'shc) : $signed(_GEN_19552); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19554 = 12'h142 == _T_643 ? $signed(7'sh15) : $signed(_GEN_19553); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19555 = 12'h143 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19554); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19556 = 12'h144 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19555); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19557 = 12'h145 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19556); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19558 = 12'h146 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19557); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19559 = 12'h147 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19558); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19560 = 12'h148 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19559); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19561 = 12'h149 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19560); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19562 = 12'h14a == _T_643 ? $signed(7'shf) : $signed(_GEN_19561); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19563 = 12'h14b == _T_643 ? $signed(7'shf) : $signed(_GEN_19562); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19564 = 12'h14c == _T_643 ? $signed(7'she) : $signed(_GEN_19563); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19565 = 12'h14d == _T_643 ? $signed(7'shd) : $signed(_GEN_19564); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19566 = 12'h14e == _T_643 ? $signed(7'shc) : $signed(_GEN_19565); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19567 = 12'h14f == _T_643 ? $signed(7'shc) : $signed(_GEN_19566); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19568 = 12'h150 == _T_643 ? $signed(7'shb) : $signed(_GEN_19567); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19569 = 12'h151 == _T_643 ? $signed(7'sha) : $signed(_GEN_19568); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19570 = 12'h152 == _T_643 ? $signed(7'sha) : $signed(_GEN_19569); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19571 = 12'h153 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19570); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19572 = 12'h154 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19571); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19573 = 12'h155 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19572); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19574 = 12'h156 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19573); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19575 = 12'h157 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19574); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19576 = 12'h158 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19575); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19577 = 12'h159 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19576); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19578 = 12'h15a == _T_643 ? $signed(7'sh4) : $signed(_GEN_19577); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19579 = 12'h15b == _T_643 ? $signed(7'sh3) : $signed(_GEN_19578); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19580 = 12'h15c == _T_643 ? $signed(7'sh3) : $signed(_GEN_19579); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19581 = 12'h15d == _T_643 ? $signed(7'sh2) : $signed(_GEN_19580); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19582 = 12'h15e == _T_643 ? $signed(7'sh1) : $signed(_GEN_19581); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19583 = 12'h15f == _T_643 ? $signed(7'sh0) : $signed(_GEN_19582); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19584 = 12'h160 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19583); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19585 = 12'h161 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19584); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19586 = 12'h162 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19585); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19587 = 12'h163 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19586); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19588 = 12'h164 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19587); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19589 = 12'h165 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19588); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19590 = 12'h166 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19589); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19591 = 12'h167 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19590); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19592 = 12'h168 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19591); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19593 = 12'h169 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19592); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19594 = 12'h16a == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19593); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19595 = 12'h16b == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19594); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19596 = 12'h16c == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19595); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19597 = 12'h16d == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19596); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19598 = 12'h16e == _T_643 ? $signed(-7'sha) : $signed(_GEN_19597); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19599 = 12'h16f == _T_643 ? $signed(-7'shb) : $signed(_GEN_19598); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19600 = 12'h170 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19599); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19601 = 12'h171 == _T_643 ? $signed(7'sh15) : $signed(_GEN_19600); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19602 = 12'h172 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19601); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19603 = 12'h173 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19602); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19604 = 12'h174 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19603); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19605 = 12'h175 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19604); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19606 = 12'h176 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19605); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19607 = 12'h177 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19606); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19608 = 12'h178 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19607); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19609 = 12'h179 == _T_643 ? $signed(7'shf) : $signed(_GEN_19608); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19610 = 12'h17a == _T_643 ? $signed(7'shf) : $signed(_GEN_19609); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19611 = 12'h17b == _T_643 ? $signed(7'she) : $signed(_GEN_19610); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19612 = 12'h17c == _T_643 ? $signed(7'shd) : $signed(_GEN_19611); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19613 = 12'h17d == _T_643 ? $signed(7'shc) : $signed(_GEN_19612); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19614 = 12'h17e == _T_643 ? $signed(7'shc) : $signed(_GEN_19613); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19615 = 12'h17f == _T_643 ? $signed(7'shb) : $signed(_GEN_19614); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19616 = 12'h180 == _T_643 ? $signed(7'sha) : $signed(_GEN_19615); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19617 = 12'h181 == _T_643 ? $signed(7'sha) : $signed(_GEN_19616); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19618 = 12'h182 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19617); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19619 = 12'h183 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19618); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19620 = 12'h184 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19619); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19621 = 12'h185 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19620); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19622 = 12'h186 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19621); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19623 = 12'h187 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19622); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19624 = 12'h188 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19623); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19625 = 12'h189 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19624); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19626 = 12'h18a == _T_643 ? $signed(7'sh3) : $signed(_GEN_19625); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19627 = 12'h18b == _T_643 ? $signed(7'sh3) : $signed(_GEN_19626); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19628 = 12'h18c == _T_643 ? $signed(7'sh2) : $signed(_GEN_19627); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19629 = 12'h18d == _T_643 ? $signed(7'sh1) : $signed(_GEN_19628); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19630 = 12'h18e == _T_643 ? $signed(7'sh0) : $signed(_GEN_19629); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19631 = 12'h18f == _T_643 ? $signed(7'sh0) : $signed(_GEN_19630); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19632 = 12'h190 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19631); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19633 = 12'h191 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19632); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19634 = 12'h192 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19633); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19635 = 12'h193 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19634); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19636 = 12'h194 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19635); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19637 = 12'h195 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19636); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19638 = 12'h196 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19637); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19639 = 12'h197 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19638); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19640 = 12'h198 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19639); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19641 = 12'h199 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19640); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19642 = 12'h19a == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19641); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19643 = 12'h19b == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19642); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19644 = 12'h19c == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19643); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19645 = 12'h19d == _T_643 ? $signed(-7'sha) : $signed(_GEN_19644); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19646 = 12'h19e == _T_643 ? $signed(7'sh16) : $signed(_GEN_19645); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19647 = 12'h19f == _T_643 ? $signed(7'sh16) : $signed(_GEN_19646); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19648 = 12'h1a0 == _T_643 ? $signed(7'sh15) : $signed(_GEN_19647); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19649 = 12'h1a1 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19648); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19650 = 12'h1a2 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19649); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19651 = 12'h1a3 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19650); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19652 = 12'h1a4 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19651); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19653 = 12'h1a5 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19652); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19654 = 12'h1a6 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19653); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19655 = 12'h1a7 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19654); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19656 = 12'h1a8 == _T_643 ? $signed(7'shf) : $signed(_GEN_19655); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19657 = 12'h1a9 == _T_643 ? $signed(7'shf) : $signed(_GEN_19656); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19658 = 12'h1aa == _T_643 ? $signed(7'she) : $signed(_GEN_19657); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19659 = 12'h1ab == _T_643 ? $signed(7'shd) : $signed(_GEN_19658); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19660 = 12'h1ac == _T_643 ? $signed(7'shc) : $signed(_GEN_19659); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19661 = 12'h1ad == _T_643 ? $signed(7'shc) : $signed(_GEN_19660); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19662 = 12'h1ae == _T_643 ? $signed(7'shb) : $signed(_GEN_19661); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19663 = 12'h1af == _T_643 ? $signed(7'sha) : $signed(_GEN_19662); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19664 = 12'h1b0 == _T_643 ? $signed(7'sha) : $signed(_GEN_19663); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19665 = 12'h1b1 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19664); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19666 = 12'h1b2 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19665); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19667 = 12'h1b3 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19666); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19668 = 12'h1b4 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19667); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19669 = 12'h1b5 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19668); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19670 = 12'h1b6 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19669); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19671 = 12'h1b7 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19670); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19672 = 12'h1b8 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19671); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19673 = 12'h1b9 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19672); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19674 = 12'h1ba == _T_643 ? $signed(7'sh3) : $signed(_GEN_19673); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19675 = 12'h1bb == _T_643 ? $signed(7'sh2) : $signed(_GEN_19674); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19676 = 12'h1bc == _T_643 ? $signed(7'sh1) : $signed(_GEN_19675); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19677 = 12'h1bd == _T_643 ? $signed(7'sh0) : $signed(_GEN_19676); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19678 = 12'h1be == _T_643 ? $signed(7'sh0) : $signed(_GEN_19677); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19679 = 12'h1bf == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19678); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19680 = 12'h1c0 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19679); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19681 = 12'h1c1 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19680); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19682 = 12'h1c2 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19681); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19683 = 12'h1c3 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19682); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19684 = 12'h1c4 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19683); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19685 = 12'h1c5 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19684); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19686 = 12'h1c6 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19685); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19687 = 12'h1c7 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19686); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19688 = 12'h1c8 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19687); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19689 = 12'h1c9 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19688); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19690 = 12'h1ca == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19689); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19691 = 12'h1cb == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19690); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19692 = 12'h1cc == _T_643 ? $signed(7'sh17) : $signed(_GEN_19691); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19693 = 12'h1cd == _T_643 ? $signed(7'sh16) : $signed(_GEN_19692); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19694 = 12'h1ce == _T_643 ? $signed(7'sh16) : $signed(_GEN_19693); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19695 = 12'h1cf == _T_643 ? $signed(7'sh15) : $signed(_GEN_19694); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19696 = 12'h1d0 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19695); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19697 = 12'h1d1 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19696); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19698 = 12'h1d2 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19697); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19699 = 12'h1d3 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19698); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19700 = 12'h1d4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19699); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19701 = 12'h1d5 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19700); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19702 = 12'h1d6 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19701); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19703 = 12'h1d7 == _T_643 ? $signed(7'shf) : $signed(_GEN_19702); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19704 = 12'h1d8 == _T_643 ? $signed(7'shf) : $signed(_GEN_19703); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19705 = 12'h1d9 == _T_643 ? $signed(7'she) : $signed(_GEN_19704); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19706 = 12'h1da == _T_643 ? $signed(7'shd) : $signed(_GEN_19705); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19707 = 12'h1db == _T_643 ? $signed(7'shc) : $signed(_GEN_19706); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19708 = 12'h1dc == _T_643 ? $signed(7'shc) : $signed(_GEN_19707); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19709 = 12'h1dd == _T_643 ? $signed(7'shb) : $signed(_GEN_19708); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19710 = 12'h1de == _T_643 ? $signed(7'sha) : $signed(_GEN_19709); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19711 = 12'h1df == _T_643 ? $signed(7'sha) : $signed(_GEN_19710); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19712 = 12'h1e0 == _T_643 ? $signed(7'sh9) : $signed(_GEN_19711); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19713 = 12'h1e1 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19712); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19714 = 12'h1e2 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19713); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19715 = 12'h1e3 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19714); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19716 = 12'h1e4 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19715); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19717 = 12'h1e5 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19716); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19718 = 12'h1e6 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19717); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19719 = 12'h1e7 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19718); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19720 = 12'h1e8 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19719); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19721 = 12'h1e9 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19720); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19722 = 12'h1ea == _T_643 ? $signed(7'sh2) : $signed(_GEN_19721); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19723 = 12'h1eb == _T_643 ? $signed(7'sh1) : $signed(_GEN_19722); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19724 = 12'h1ec == _T_643 ? $signed(7'sh0) : $signed(_GEN_19723); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19725 = 12'h1ed == _T_643 ? $signed(7'sh0) : $signed(_GEN_19724); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19726 = 12'h1ee == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19725); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19727 = 12'h1ef == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19726); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19728 = 12'h1f0 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19727); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19729 = 12'h1f1 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19728); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19730 = 12'h1f2 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19729); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19731 = 12'h1f3 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19730); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19732 = 12'h1f4 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19731); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19733 = 12'h1f5 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19732); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19734 = 12'h1f6 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19733); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19735 = 12'h1f7 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19734); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19736 = 12'h1f8 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19735); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19737 = 12'h1f9 == _T_643 ? $signed(-7'sh9) : $signed(_GEN_19736); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19738 = 12'h1fa == _T_643 ? $signed(7'sh18) : $signed(_GEN_19737); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19739 = 12'h1fb == _T_643 ? $signed(7'sh17) : $signed(_GEN_19738); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19740 = 12'h1fc == _T_643 ? $signed(7'sh16) : $signed(_GEN_19739); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19741 = 12'h1fd == _T_643 ? $signed(7'sh16) : $signed(_GEN_19740); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19742 = 12'h1fe == _T_643 ? $signed(7'sh15) : $signed(_GEN_19741); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19743 = 12'h1ff == _T_643 ? $signed(7'sh14) : $signed(_GEN_19742); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19744 = 12'h200 == _T_643 ? $signed(7'sh14) : $signed(_GEN_19743); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19745 = 12'h201 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19744); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19746 = 12'h202 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19745); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19747 = 12'h203 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19746); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19748 = 12'h204 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19747); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19749 = 12'h205 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19748); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19750 = 12'h206 == _T_643 ? $signed(7'shf) : $signed(_GEN_19749); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19751 = 12'h207 == _T_643 ? $signed(7'shf) : $signed(_GEN_19750); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19752 = 12'h208 == _T_643 ? $signed(7'she) : $signed(_GEN_19751); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19753 = 12'h209 == _T_643 ? $signed(7'shd) : $signed(_GEN_19752); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19754 = 12'h20a == _T_643 ? $signed(7'shc) : $signed(_GEN_19753); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19755 = 12'h20b == _T_643 ? $signed(7'shc) : $signed(_GEN_19754); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19756 = 12'h20c == _T_643 ? $signed(7'shb) : $signed(_GEN_19755); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19757 = 12'h20d == _T_643 ? $signed(7'sha) : $signed(_GEN_19756); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19758 = 12'h20e == _T_643 ? $signed(7'sha) : $signed(_GEN_19757); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19759 = 12'h20f == _T_643 ? $signed(7'sh9) : $signed(_GEN_19758); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19760 = 12'h210 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19759); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19761 = 12'h211 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19760); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19762 = 12'h212 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19761); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19763 = 12'h213 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19762); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19764 = 12'h214 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19763); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19765 = 12'h215 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19764); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19766 = 12'h216 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19765); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19767 = 12'h217 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19766); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19768 = 12'h218 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19767); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19769 = 12'h219 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19768); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19770 = 12'h21a == _T_643 ? $signed(7'sh1) : $signed(_GEN_19769); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19771 = 12'h21b == _T_643 ? $signed(7'sh0) : $signed(_GEN_19770); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19772 = 12'h21c == _T_643 ? $signed(7'sh0) : $signed(_GEN_19771); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19773 = 12'h21d == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19772); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19774 = 12'h21e == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19773); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19775 = 12'h21f == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19774); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19776 = 12'h220 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19775); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19777 = 12'h221 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19776); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19778 = 12'h222 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19777); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19779 = 12'h223 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19778); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19780 = 12'h224 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19779); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19781 = 12'h225 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19780); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19782 = 12'h226 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19781); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19783 = 12'h227 == _T_643 ? $signed(-7'sh8) : $signed(_GEN_19782); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19784 = 12'h228 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19783); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19785 = 12'h229 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19784); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19786 = 12'h22a == _T_643 ? $signed(7'sh17) : $signed(_GEN_19785); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19787 = 12'h22b == _T_643 ? $signed(7'sh16) : $signed(_GEN_19786); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19788 = 12'h22c == _T_643 ? $signed(7'sh16) : $signed(_GEN_19787); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19789 = 12'h22d == _T_643 ? $signed(7'sh15) : $signed(_GEN_19788); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19790 = 12'h22e == _T_643 ? $signed(7'sh14) : $signed(_GEN_19789); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19791 = 12'h22f == _T_643 ? $signed(7'sh14) : $signed(_GEN_19790); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19792 = 12'h230 == _T_643 ? $signed(7'sh13) : $signed(_GEN_19791); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19793 = 12'h231 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19792); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19794 = 12'h232 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19793); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19795 = 12'h233 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19794); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19796 = 12'h234 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19795); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19797 = 12'h235 == _T_643 ? $signed(7'shf) : $signed(_GEN_19796); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19798 = 12'h236 == _T_643 ? $signed(7'shf) : $signed(_GEN_19797); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19799 = 12'h237 == _T_643 ? $signed(7'she) : $signed(_GEN_19798); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19800 = 12'h238 == _T_643 ? $signed(7'shd) : $signed(_GEN_19799); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19801 = 12'h239 == _T_643 ? $signed(7'shc) : $signed(_GEN_19800); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19802 = 12'h23a == _T_643 ? $signed(7'shc) : $signed(_GEN_19801); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19803 = 12'h23b == _T_643 ? $signed(7'shb) : $signed(_GEN_19802); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19804 = 12'h23c == _T_643 ? $signed(7'sha) : $signed(_GEN_19803); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19805 = 12'h23d == _T_643 ? $signed(7'sha) : $signed(_GEN_19804); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19806 = 12'h23e == _T_643 ? $signed(7'sh9) : $signed(_GEN_19805); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19807 = 12'h23f == _T_643 ? $signed(7'sh8) : $signed(_GEN_19806); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19808 = 12'h240 == _T_643 ? $signed(7'sh8) : $signed(_GEN_19807); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19809 = 12'h241 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19808); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19810 = 12'h242 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19809); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19811 = 12'h243 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19810); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19812 = 12'h244 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19811); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19813 = 12'h245 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19812); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19814 = 12'h246 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19813); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19815 = 12'h247 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19814); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19816 = 12'h248 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19815); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19817 = 12'h249 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19816); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19818 = 12'h24a == _T_643 ? $signed(7'sh0) : $signed(_GEN_19817); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19819 = 12'h24b == _T_643 ? $signed(7'sh0) : $signed(_GEN_19818); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19820 = 12'h24c == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19819); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19821 = 12'h24d == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19820); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19822 = 12'h24e == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19821); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19823 = 12'h24f == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19822); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19824 = 12'h250 == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19823); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19825 = 12'h251 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19824); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19826 = 12'h252 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19825); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19827 = 12'h253 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19826); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19828 = 12'h254 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19827); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19829 = 12'h255 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19828); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19830 = 12'h256 == _T_643 ? $signed(7'sh19) : $signed(_GEN_19829); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19831 = 12'h257 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19830); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19832 = 12'h258 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19831); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19833 = 12'h259 == _T_643 ? $signed(7'sh17) : $signed(_GEN_19832); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19834 = 12'h25a == _T_643 ? $signed(7'sh16) : $signed(_GEN_19833); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19835 = 12'h25b == _T_643 ? $signed(7'sh16) : $signed(_GEN_19834); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19836 = 12'h25c == _T_643 ? $signed(7'sh15) : $signed(_GEN_19835); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19837 = 12'h25d == _T_643 ? $signed(7'sh14) : $signed(_GEN_19836); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19838 = 12'h25e == _T_643 ? $signed(7'sh14) : $signed(_GEN_19837); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19839 = 12'h25f == _T_643 ? $signed(7'sh13) : $signed(_GEN_19838); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19840 = 12'h260 == _T_643 ? $signed(7'sh12) : $signed(_GEN_19839); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19841 = 12'h261 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19840); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19842 = 12'h262 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19841); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19843 = 12'h263 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19842); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19844 = 12'h264 == _T_643 ? $signed(7'shf) : $signed(_GEN_19843); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19845 = 12'h265 == _T_643 ? $signed(7'shf) : $signed(_GEN_19844); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19846 = 12'h266 == _T_643 ? $signed(7'she) : $signed(_GEN_19845); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19847 = 12'h267 == _T_643 ? $signed(7'shd) : $signed(_GEN_19846); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19848 = 12'h268 == _T_643 ? $signed(7'shc) : $signed(_GEN_19847); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19849 = 12'h269 == _T_643 ? $signed(7'shc) : $signed(_GEN_19848); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19850 = 12'h26a == _T_643 ? $signed(7'shb) : $signed(_GEN_19849); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19851 = 12'h26b == _T_643 ? $signed(7'sha) : $signed(_GEN_19850); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19852 = 12'h26c == _T_643 ? $signed(7'sha) : $signed(_GEN_19851); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19853 = 12'h26d == _T_643 ? $signed(7'sh9) : $signed(_GEN_19852); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19854 = 12'h26e == _T_643 ? $signed(7'sh8) : $signed(_GEN_19853); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19855 = 12'h26f == _T_643 ? $signed(7'sh8) : $signed(_GEN_19854); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19856 = 12'h270 == _T_643 ? $signed(7'sh7) : $signed(_GEN_19855); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19857 = 12'h271 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19856); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19858 = 12'h272 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19857); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19859 = 12'h273 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19858); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19860 = 12'h274 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19859); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19861 = 12'h275 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19860); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19862 = 12'h276 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19861); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19863 = 12'h277 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19862); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19864 = 12'h278 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19863); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19865 = 12'h279 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19864); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19866 = 12'h27a == _T_643 ? $signed(7'sh0) : $signed(_GEN_19865); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19867 = 12'h27b == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19866); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19868 = 12'h27c == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19867); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19869 = 12'h27d == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19868); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19870 = 12'h27e == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19869); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19871 = 12'h27f == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19870); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19872 = 12'h280 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19871); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19873 = 12'h281 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19872); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19874 = 12'h282 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19873); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19875 = 12'h283 == _T_643 ? $signed(-7'sh7) : $signed(_GEN_19874); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19876 = 12'h284 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19875); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19877 = 12'h285 == _T_643 ? $signed(7'sh19) : $signed(_GEN_19876); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19878 = 12'h286 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19877); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19879 = 12'h287 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19878); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19880 = 12'h288 == _T_643 ? $signed(7'sh17) : $signed(_GEN_19879); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19881 = 12'h289 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19880); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19882 = 12'h28a == _T_643 ? $signed(7'sh16) : $signed(_GEN_19881); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19883 = 12'h28b == _T_643 ? $signed(7'sh15) : $signed(_GEN_19882); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19884 = 12'h28c == _T_643 ? $signed(7'sh14) : $signed(_GEN_19883); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19885 = 12'h28d == _T_643 ? $signed(7'sh14) : $signed(_GEN_19884); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19886 = 12'h28e == _T_643 ? $signed(7'sh13) : $signed(_GEN_19885); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19887 = 12'h28f == _T_643 ? $signed(7'sh12) : $signed(_GEN_19886); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19888 = 12'h290 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19887); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19889 = 12'h291 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19888); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19890 = 12'h292 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19889); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19891 = 12'h293 == _T_643 ? $signed(7'shf) : $signed(_GEN_19890); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19892 = 12'h294 == _T_643 ? $signed(7'shf) : $signed(_GEN_19891); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19893 = 12'h295 == _T_643 ? $signed(7'she) : $signed(_GEN_19892); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19894 = 12'h296 == _T_643 ? $signed(7'shd) : $signed(_GEN_19893); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19895 = 12'h297 == _T_643 ? $signed(7'shc) : $signed(_GEN_19894); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19896 = 12'h298 == _T_643 ? $signed(7'shc) : $signed(_GEN_19895); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19897 = 12'h299 == _T_643 ? $signed(7'shb) : $signed(_GEN_19896); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19898 = 12'h29a == _T_643 ? $signed(7'sha) : $signed(_GEN_19897); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19899 = 12'h29b == _T_643 ? $signed(7'sha) : $signed(_GEN_19898); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19900 = 12'h29c == _T_643 ? $signed(7'sh9) : $signed(_GEN_19899); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19901 = 12'h29d == _T_643 ? $signed(7'sh8) : $signed(_GEN_19900); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19902 = 12'h29e == _T_643 ? $signed(7'sh8) : $signed(_GEN_19901); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19903 = 12'h29f == _T_643 ? $signed(7'sh7) : $signed(_GEN_19902); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19904 = 12'h2a0 == _T_643 ? $signed(7'sh6) : $signed(_GEN_19903); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19905 = 12'h2a1 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19904); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19906 = 12'h2a2 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19905); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19907 = 12'h2a3 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19906); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19908 = 12'h2a4 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19907); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19909 = 12'h2a5 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19908); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19910 = 12'h2a6 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19909); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19911 = 12'h2a7 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19910); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19912 = 12'h2a8 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19911); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19913 = 12'h2a9 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19912); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19914 = 12'h2aa == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19913); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19915 = 12'h2ab == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19914); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19916 = 12'h2ac == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19915); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19917 = 12'h2ad == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19916); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19918 = 12'h2ae == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19917); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19919 = 12'h2af == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19918); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19920 = 12'h2b0 == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19919); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19921 = 12'h2b1 == _T_643 ? $signed(-7'sh6) : $signed(_GEN_19920); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19922 = 12'h2b2 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19921); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19923 = 12'h2b3 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19922); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19924 = 12'h2b4 == _T_643 ? $signed(7'sh19) : $signed(_GEN_19923); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19925 = 12'h2b5 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19924); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19926 = 12'h2b6 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19925); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19927 = 12'h2b7 == _T_643 ? $signed(7'sh17) : $signed(_GEN_19926); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19928 = 12'h2b8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19927); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19929 = 12'h2b9 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19928); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19930 = 12'h2ba == _T_643 ? $signed(7'sh15) : $signed(_GEN_19929); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19931 = 12'h2bb == _T_643 ? $signed(7'sh14) : $signed(_GEN_19930); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19932 = 12'h2bc == _T_643 ? $signed(7'sh14) : $signed(_GEN_19931); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19933 = 12'h2bd == _T_643 ? $signed(7'sh13) : $signed(_GEN_19932); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19934 = 12'h2be == _T_643 ? $signed(7'sh12) : $signed(_GEN_19933); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19935 = 12'h2bf == _T_643 ? $signed(7'sh11) : $signed(_GEN_19934); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19936 = 12'h2c0 == _T_643 ? $signed(7'sh11) : $signed(_GEN_19935); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19937 = 12'h2c1 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19936); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19938 = 12'h2c2 == _T_643 ? $signed(7'shf) : $signed(_GEN_19937); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19939 = 12'h2c3 == _T_643 ? $signed(7'shf) : $signed(_GEN_19938); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19940 = 12'h2c4 == _T_643 ? $signed(7'she) : $signed(_GEN_19939); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19941 = 12'h2c5 == _T_643 ? $signed(7'shd) : $signed(_GEN_19940); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19942 = 12'h2c6 == _T_643 ? $signed(7'shc) : $signed(_GEN_19941); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19943 = 12'h2c7 == _T_643 ? $signed(7'shc) : $signed(_GEN_19942); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19944 = 12'h2c8 == _T_643 ? $signed(7'shb) : $signed(_GEN_19943); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19945 = 12'h2c9 == _T_643 ? $signed(7'sha) : $signed(_GEN_19944); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19946 = 12'h2ca == _T_643 ? $signed(7'sha) : $signed(_GEN_19945); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19947 = 12'h2cb == _T_643 ? $signed(7'sh9) : $signed(_GEN_19946); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19948 = 12'h2cc == _T_643 ? $signed(7'sh8) : $signed(_GEN_19947); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19949 = 12'h2cd == _T_643 ? $signed(7'sh8) : $signed(_GEN_19948); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19950 = 12'h2ce == _T_643 ? $signed(7'sh7) : $signed(_GEN_19949); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19951 = 12'h2cf == _T_643 ? $signed(7'sh6) : $signed(_GEN_19950); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19952 = 12'h2d0 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19951); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19953 = 12'h2d1 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19952); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19954 = 12'h2d2 == _T_643 ? $signed(7'sh4) : $signed(_GEN_19953); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19955 = 12'h2d3 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19954); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19956 = 12'h2d4 == _T_643 ? $signed(7'sh3) : $signed(_GEN_19955); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19957 = 12'h2d5 == _T_643 ? $signed(7'sh2) : $signed(_GEN_19956); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19958 = 12'h2d6 == _T_643 ? $signed(7'sh1) : $signed(_GEN_19957); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19959 = 12'h2d7 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19958); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19960 = 12'h2d8 == _T_643 ? $signed(7'sh0) : $signed(_GEN_19959); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19961 = 12'h2d9 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_19960); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19962 = 12'h2da == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19961); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19963 = 12'h2db == _T_643 ? $signed(-7'sh2) : $signed(_GEN_19962); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19964 = 12'h2dc == _T_643 ? $signed(-7'sh3) : $signed(_GEN_19963); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19965 = 12'h2dd == _T_643 ? $signed(-7'sh4) : $signed(_GEN_19964); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19966 = 12'h2de == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19965); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19967 = 12'h2df == _T_643 ? $signed(-7'sh5) : $signed(_GEN_19966); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19968 = 12'h2e0 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19967); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19969 = 12'h2e1 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_19968); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19970 = 12'h2e2 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_19969); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19971 = 12'h2e3 == _T_643 ? $signed(7'sh19) : $signed(_GEN_19970); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19972 = 12'h2e4 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19971); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19973 = 12'h2e5 == _T_643 ? $signed(7'sh18) : $signed(_GEN_19972); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19974 = 12'h2e6 == _T_643 ? $signed(7'sh17) : $signed(_GEN_19973); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19975 = 12'h2e7 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19974); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19976 = 12'h2e8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_19975); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19977 = 12'h2e9 == _T_643 ? $signed(7'sh15) : $signed(_GEN_19976); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19978 = 12'h2ea == _T_643 ? $signed(7'sh14) : $signed(_GEN_19977); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19979 = 12'h2eb == _T_643 ? $signed(7'sh14) : $signed(_GEN_19978); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19980 = 12'h2ec == _T_643 ? $signed(7'sh13) : $signed(_GEN_19979); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19981 = 12'h2ed == _T_643 ? $signed(7'sh12) : $signed(_GEN_19980); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19982 = 12'h2ee == _T_643 ? $signed(7'sh11) : $signed(_GEN_19981); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19983 = 12'h2ef == _T_643 ? $signed(7'sh11) : $signed(_GEN_19982); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19984 = 12'h2f0 == _T_643 ? $signed(7'sh10) : $signed(_GEN_19983); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19985 = 12'h2f1 == _T_643 ? $signed(7'shf) : $signed(_GEN_19984); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19986 = 12'h2f2 == _T_643 ? $signed(7'shf) : $signed(_GEN_19985); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19987 = 12'h2f3 == _T_643 ? $signed(7'she) : $signed(_GEN_19986); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19988 = 12'h2f4 == _T_643 ? $signed(7'shd) : $signed(_GEN_19987); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19989 = 12'h2f5 == _T_643 ? $signed(7'shc) : $signed(_GEN_19988); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19990 = 12'h2f6 == _T_643 ? $signed(7'shc) : $signed(_GEN_19989); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19991 = 12'h2f7 == _T_643 ? $signed(7'shb) : $signed(_GEN_19990); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19992 = 12'h2f8 == _T_643 ? $signed(7'sha) : $signed(_GEN_19991); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19993 = 12'h2f9 == _T_643 ? $signed(7'sha) : $signed(_GEN_19992); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19994 = 12'h2fa == _T_643 ? $signed(7'sh9) : $signed(_GEN_19993); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19995 = 12'h2fb == _T_643 ? $signed(7'sh8) : $signed(_GEN_19994); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19996 = 12'h2fc == _T_643 ? $signed(7'sh8) : $signed(_GEN_19995); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19997 = 12'h2fd == _T_643 ? $signed(7'sh7) : $signed(_GEN_19996); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19998 = 12'h2fe == _T_643 ? $signed(7'sh6) : $signed(_GEN_19997); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_19999 = 12'h2ff == _T_643 ? $signed(7'sh5) : $signed(_GEN_19998); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20000 = 12'h300 == _T_643 ? $signed(7'sh5) : $signed(_GEN_19999); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20001 = 12'h301 == _T_643 ? $signed(7'sh4) : $signed(_GEN_20000); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20002 = 12'h302 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20001); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20003 = 12'h303 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20002); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20004 = 12'h304 == _T_643 ? $signed(7'sh2) : $signed(_GEN_20003); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20005 = 12'h305 == _T_643 ? $signed(7'sh1) : $signed(_GEN_20004); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20006 = 12'h306 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20005); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20007 = 12'h307 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20006); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20008 = 12'h308 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_20007); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20009 = 12'h309 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20008); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20010 = 12'h30a == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20009); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20011 = 12'h30b == _T_643 ? $signed(-7'sh3) : $signed(_GEN_20010); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20012 = 12'h30c == _T_643 ? $signed(-7'sh4) : $signed(_GEN_20011); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20013 = 12'h30d == _T_643 ? $signed(-7'sh5) : $signed(_GEN_20012); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20014 = 12'h30e == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20013); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20015 = 12'h30f == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20014); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20016 = 12'h310 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20015); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20017 = 12'h311 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20016); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20018 = 12'h312 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20017); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20019 = 12'h313 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20018); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20020 = 12'h314 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20019); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20021 = 12'h315 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20020); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20022 = 12'h316 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20021); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20023 = 12'h317 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20022); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20024 = 12'h318 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20023); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20025 = 12'h319 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20024); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20026 = 12'h31a == _T_643 ? $signed(7'sh14) : $signed(_GEN_20025); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20027 = 12'h31b == _T_643 ? $signed(7'sh13) : $signed(_GEN_20026); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20028 = 12'h31c == _T_643 ? $signed(7'sh12) : $signed(_GEN_20027); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20029 = 12'h31d == _T_643 ? $signed(7'sh11) : $signed(_GEN_20028); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20030 = 12'h31e == _T_643 ? $signed(7'sh11) : $signed(_GEN_20029); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20031 = 12'h31f == _T_643 ? $signed(7'sh10) : $signed(_GEN_20030); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20032 = 12'h320 == _T_643 ? $signed(7'shf) : $signed(_GEN_20031); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20033 = 12'h321 == _T_643 ? $signed(7'shf) : $signed(_GEN_20032); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20034 = 12'h322 == _T_643 ? $signed(7'she) : $signed(_GEN_20033); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20035 = 12'h323 == _T_643 ? $signed(7'shd) : $signed(_GEN_20034); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20036 = 12'h324 == _T_643 ? $signed(7'shc) : $signed(_GEN_20035); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20037 = 12'h325 == _T_643 ? $signed(7'shc) : $signed(_GEN_20036); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20038 = 12'h326 == _T_643 ? $signed(7'shb) : $signed(_GEN_20037); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20039 = 12'h327 == _T_643 ? $signed(7'sha) : $signed(_GEN_20038); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20040 = 12'h328 == _T_643 ? $signed(7'sha) : $signed(_GEN_20039); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20041 = 12'h329 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20040); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20042 = 12'h32a == _T_643 ? $signed(7'sh8) : $signed(_GEN_20041); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20043 = 12'h32b == _T_643 ? $signed(7'sh8) : $signed(_GEN_20042); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20044 = 12'h32c == _T_643 ? $signed(7'sh7) : $signed(_GEN_20043); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20045 = 12'h32d == _T_643 ? $signed(7'sh6) : $signed(_GEN_20044); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20046 = 12'h32e == _T_643 ? $signed(7'sh5) : $signed(_GEN_20045); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20047 = 12'h32f == _T_643 ? $signed(7'sh5) : $signed(_GEN_20046); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20048 = 12'h330 == _T_643 ? $signed(7'sh4) : $signed(_GEN_20047); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20049 = 12'h331 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20048); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20050 = 12'h332 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20049); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20051 = 12'h333 == _T_643 ? $signed(7'sh2) : $signed(_GEN_20050); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20052 = 12'h334 == _T_643 ? $signed(7'sh1) : $signed(_GEN_20051); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20053 = 12'h335 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20052); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20054 = 12'h336 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20053); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20055 = 12'h337 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_20054); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20056 = 12'h338 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20055); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20057 = 12'h339 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20056); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20058 = 12'h33a == _T_643 ? $signed(-7'sh3) : $signed(_GEN_20057); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20059 = 12'h33b == _T_643 ? $signed(-7'sh4) : $signed(_GEN_20058); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20060 = 12'h33c == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20059); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20061 = 12'h33d == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20060); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20062 = 12'h33e == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20061); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20063 = 12'h33f == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20062); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20064 = 12'h340 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20063); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20065 = 12'h341 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20064); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20066 = 12'h342 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20065); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20067 = 12'h343 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20066); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20068 = 12'h344 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20067); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20069 = 12'h345 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20068); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20070 = 12'h346 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20069); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20071 = 12'h347 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20070); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20072 = 12'h348 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20071); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20073 = 12'h349 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20072); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20074 = 12'h34a == _T_643 ? $signed(7'sh13) : $signed(_GEN_20073); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20075 = 12'h34b == _T_643 ? $signed(7'sh12) : $signed(_GEN_20074); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20076 = 12'h34c == _T_643 ? $signed(7'sh11) : $signed(_GEN_20075); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20077 = 12'h34d == _T_643 ? $signed(7'sh11) : $signed(_GEN_20076); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20078 = 12'h34e == _T_643 ? $signed(7'sh10) : $signed(_GEN_20077); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20079 = 12'h34f == _T_643 ? $signed(7'shf) : $signed(_GEN_20078); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20080 = 12'h350 == _T_643 ? $signed(7'shf) : $signed(_GEN_20079); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20081 = 12'h351 == _T_643 ? $signed(7'she) : $signed(_GEN_20080); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20082 = 12'h352 == _T_643 ? $signed(7'shd) : $signed(_GEN_20081); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20083 = 12'h353 == _T_643 ? $signed(7'shc) : $signed(_GEN_20082); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20084 = 12'h354 == _T_643 ? $signed(7'shc) : $signed(_GEN_20083); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20085 = 12'h355 == _T_643 ? $signed(7'shb) : $signed(_GEN_20084); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20086 = 12'h356 == _T_643 ? $signed(7'sha) : $signed(_GEN_20085); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20087 = 12'h357 == _T_643 ? $signed(7'sha) : $signed(_GEN_20086); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20088 = 12'h358 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20087); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20089 = 12'h359 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20088); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20090 = 12'h35a == _T_643 ? $signed(7'sh8) : $signed(_GEN_20089); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20091 = 12'h35b == _T_643 ? $signed(7'sh7) : $signed(_GEN_20090); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20092 = 12'h35c == _T_643 ? $signed(7'sh6) : $signed(_GEN_20091); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20093 = 12'h35d == _T_643 ? $signed(7'sh5) : $signed(_GEN_20092); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20094 = 12'h35e == _T_643 ? $signed(7'sh5) : $signed(_GEN_20093); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20095 = 12'h35f == _T_643 ? $signed(7'sh4) : $signed(_GEN_20094); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20096 = 12'h360 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20095); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20097 = 12'h361 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20096); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20098 = 12'h362 == _T_643 ? $signed(7'sh2) : $signed(_GEN_20097); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20099 = 12'h363 == _T_643 ? $signed(7'sh1) : $signed(_GEN_20098); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20100 = 12'h364 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20099); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20101 = 12'h365 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20100); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20102 = 12'h366 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_20101); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20103 = 12'h367 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20102); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20104 = 12'h368 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20103); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20105 = 12'h369 == _T_643 ? $signed(-7'sh3) : $signed(_GEN_20104); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20106 = 12'h36a == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20105); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20107 = 12'h36b == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20106); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20108 = 12'h36c == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20107); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20109 = 12'h36d == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20108); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20110 = 12'h36e == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20109); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20111 = 12'h36f == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20110); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20112 = 12'h370 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20111); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20113 = 12'h371 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20112); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20114 = 12'h372 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20113); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20115 = 12'h373 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20114); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20116 = 12'h374 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20115); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20117 = 12'h375 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20116); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20118 = 12'h376 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20117); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20119 = 12'h377 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20118); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20120 = 12'h378 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20119); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20121 = 12'h379 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20120); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20122 = 12'h37a == _T_643 ? $signed(7'sh12) : $signed(_GEN_20121); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20123 = 12'h37b == _T_643 ? $signed(7'sh11) : $signed(_GEN_20122); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20124 = 12'h37c == _T_643 ? $signed(7'sh11) : $signed(_GEN_20123); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20125 = 12'h37d == _T_643 ? $signed(7'sh10) : $signed(_GEN_20124); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20126 = 12'h37e == _T_643 ? $signed(7'shf) : $signed(_GEN_20125); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20127 = 12'h37f == _T_643 ? $signed(7'shf) : $signed(_GEN_20126); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20128 = 12'h380 == _T_643 ? $signed(7'she) : $signed(_GEN_20127); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20129 = 12'h381 == _T_643 ? $signed(7'shd) : $signed(_GEN_20128); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20130 = 12'h382 == _T_643 ? $signed(7'shc) : $signed(_GEN_20129); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20131 = 12'h383 == _T_643 ? $signed(7'shc) : $signed(_GEN_20130); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20132 = 12'h384 == _T_643 ? $signed(7'shb) : $signed(_GEN_20131); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20133 = 12'h385 == _T_643 ? $signed(7'sha) : $signed(_GEN_20132); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20134 = 12'h386 == _T_643 ? $signed(7'sha) : $signed(_GEN_20133); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20135 = 12'h387 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20134); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20136 = 12'h388 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20135); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20137 = 12'h389 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20136); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20138 = 12'h38a == _T_643 ? $signed(7'sh7) : $signed(_GEN_20137); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20139 = 12'h38b == _T_643 ? $signed(7'sh6) : $signed(_GEN_20138); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20140 = 12'h38c == _T_643 ? $signed(7'sh5) : $signed(_GEN_20139); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20141 = 12'h38d == _T_643 ? $signed(7'sh5) : $signed(_GEN_20140); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20142 = 12'h38e == _T_643 ? $signed(7'sh4) : $signed(_GEN_20141); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20143 = 12'h38f == _T_643 ? $signed(7'sh3) : $signed(_GEN_20142); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20144 = 12'h390 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20143); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20145 = 12'h391 == _T_643 ? $signed(7'sh2) : $signed(_GEN_20144); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20146 = 12'h392 == _T_643 ? $signed(7'sh1) : $signed(_GEN_20145); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20147 = 12'h393 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20146); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20148 = 12'h394 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20147); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20149 = 12'h395 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_20148); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20150 = 12'h396 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20149); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20151 = 12'h397 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20150); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20152 = 12'h398 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20151); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20153 = 12'h399 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20152); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20154 = 12'h39a == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20153); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20155 = 12'h39b == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20154); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20156 = 12'h39c == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20155); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20157 = 12'h39d == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20156); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20158 = 12'h39e == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20157); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20159 = 12'h39f == _T_643 ? $signed(7'sh19) : $signed(_GEN_20158); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20160 = 12'h3a0 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20159); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20161 = 12'h3a1 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20160); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20162 = 12'h3a2 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20161); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20163 = 12'h3a3 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20162); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20164 = 12'h3a4 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20163); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20165 = 12'h3a5 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20164); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20166 = 12'h3a6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20165); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20167 = 12'h3a7 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20166); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20168 = 12'h3a8 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20167); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20169 = 12'h3a9 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20168); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20170 = 12'h3aa == _T_643 ? $signed(7'sh11) : $signed(_GEN_20169); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20171 = 12'h3ab == _T_643 ? $signed(7'sh11) : $signed(_GEN_20170); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20172 = 12'h3ac == _T_643 ? $signed(7'sh10) : $signed(_GEN_20171); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20173 = 12'h3ad == _T_643 ? $signed(7'shf) : $signed(_GEN_20172); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20174 = 12'h3ae == _T_643 ? $signed(7'shf) : $signed(_GEN_20173); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20175 = 12'h3af == _T_643 ? $signed(7'she) : $signed(_GEN_20174); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20176 = 12'h3b0 == _T_643 ? $signed(7'shd) : $signed(_GEN_20175); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20177 = 12'h3b1 == _T_643 ? $signed(7'shc) : $signed(_GEN_20176); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20178 = 12'h3b2 == _T_643 ? $signed(7'shc) : $signed(_GEN_20177); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20179 = 12'h3b3 == _T_643 ? $signed(7'shb) : $signed(_GEN_20178); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20180 = 12'h3b4 == _T_643 ? $signed(7'sha) : $signed(_GEN_20179); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20181 = 12'h3b5 == _T_643 ? $signed(7'sha) : $signed(_GEN_20180); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20182 = 12'h3b6 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20181); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20183 = 12'h3b7 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20182); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20184 = 12'h3b8 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20183); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20185 = 12'h3b9 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20184); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20186 = 12'h3ba == _T_643 ? $signed(7'sh6) : $signed(_GEN_20185); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20187 = 12'h3bb == _T_643 ? $signed(7'sh5) : $signed(_GEN_20186); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20188 = 12'h3bc == _T_643 ? $signed(7'sh5) : $signed(_GEN_20187); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20189 = 12'h3bd == _T_643 ? $signed(7'sh4) : $signed(_GEN_20188); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20190 = 12'h3be == _T_643 ? $signed(7'sh3) : $signed(_GEN_20189); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20191 = 12'h3bf == _T_643 ? $signed(7'sh3) : $signed(_GEN_20190); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20192 = 12'h3c0 == _T_643 ? $signed(7'sh2) : $signed(_GEN_20191); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20193 = 12'h3c1 == _T_643 ? $signed(7'sh1) : $signed(_GEN_20192); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20194 = 12'h3c2 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20193); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20195 = 12'h3c3 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20194); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20196 = 12'h3c4 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_20195); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20197 = 12'h3c5 == _T_643 ? $signed(-7'sh2) : $signed(_GEN_20196); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20198 = 12'h3c6 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20197); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20199 = 12'h3c7 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20198); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20200 = 12'h3c8 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20199); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20201 = 12'h3c9 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20200); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20202 = 12'h3ca == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20201); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20203 = 12'h3cb == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20202); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20204 = 12'h3cc == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20203); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20205 = 12'h3cd == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20204); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20206 = 12'h3ce == _T_643 ? $signed(7'sh19) : $signed(_GEN_20205); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20207 = 12'h3cf == _T_643 ? $signed(7'sh18) : $signed(_GEN_20206); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20208 = 12'h3d0 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20207); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20209 = 12'h3d1 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20208); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20210 = 12'h3d2 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20209); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20211 = 12'h3d3 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20210); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20212 = 12'h3d4 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20211); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20213 = 12'h3d5 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20212); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20214 = 12'h3d6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20213); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20215 = 12'h3d7 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20214); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20216 = 12'h3d8 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20215); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20217 = 12'h3d9 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20216); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20218 = 12'h3da == _T_643 ? $signed(7'sh11) : $signed(_GEN_20217); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20219 = 12'h3db == _T_643 ? $signed(7'sh10) : $signed(_GEN_20218); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20220 = 12'h3dc == _T_643 ? $signed(7'shf) : $signed(_GEN_20219); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20221 = 12'h3dd == _T_643 ? $signed(7'shf) : $signed(_GEN_20220); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20222 = 12'h3de == _T_643 ? $signed(7'she) : $signed(_GEN_20221); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20223 = 12'h3df == _T_643 ? $signed(7'shd) : $signed(_GEN_20222); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20224 = 12'h3e0 == _T_643 ? $signed(7'shc) : $signed(_GEN_20223); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20225 = 12'h3e1 == _T_643 ? $signed(7'shc) : $signed(_GEN_20224); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20226 = 12'h3e2 == _T_643 ? $signed(7'shb) : $signed(_GEN_20225); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20227 = 12'h3e3 == _T_643 ? $signed(7'sha) : $signed(_GEN_20226); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20228 = 12'h3e4 == _T_643 ? $signed(7'sha) : $signed(_GEN_20227); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20229 = 12'h3e5 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20228); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20230 = 12'h3e6 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20229); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20231 = 12'h3e7 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20230); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20232 = 12'h3e8 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20231); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20233 = 12'h3e9 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20232); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20234 = 12'h3ea == _T_643 ? $signed(7'sh5) : $signed(_GEN_20233); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20235 = 12'h3eb == _T_643 ? $signed(7'sh5) : $signed(_GEN_20234); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20236 = 12'h3ec == _T_643 ? $signed(7'sh4) : $signed(_GEN_20235); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20237 = 12'h3ed == _T_643 ? $signed(7'sh3) : $signed(_GEN_20236); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20238 = 12'h3ee == _T_643 ? $signed(7'sh3) : $signed(_GEN_20237); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20239 = 12'h3ef == _T_643 ? $signed(7'sh2) : $signed(_GEN_20238); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20240 = 12'h3f0 == _T_643 ? $signed(7'sh1) : $signed(_GEN_20239); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20241 = 12'h3f1 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20240); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20242 = 12'h3f2 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20241); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20243 = 12'h3f3 == _T_643 ? $signed(-7'sh1) : $signed(_GEN_20242); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20244 = 12'h3f4 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20243); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20245 = 12'h3f5 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20244); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20246 = 12'h3f6 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20245); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20247 = 12'h3f7 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20246); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20248 = 12'h3f8 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20247); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20249 = 12'h3f9 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20248); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20250 = 12'h3fa == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20249); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20251 = 12'h3fb == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20250); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20252 = 12'h3fc == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20251); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20253 = 12'h3fd == _T_643 ? $signed(7'sh19) : $signed(_GEN_20252); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20254 = 12'h3fe == _T_643 ? $signed(7'sh18) : $signed(_GEN_20253); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20255 = 12'h3ff == _T_643 ? $signed(7'sh18) : $signed(_GEN_20254); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20256 = 12'h400 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20255); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20257 = 12'h401 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20256); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20258 = 12'h402 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20257); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20259 = 12'h403 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20258); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20260 = 12'h404 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20259); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20261 = 12'h405 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20260); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20262 = 12'h406 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20261); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20263 = 12'h407 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20262); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20264 = 12'h408 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20263); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20265 = 12'h409 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20264); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20266 = 12'h40a == _T_643 ? $signed(7'sh10) : $signed(_GEN_20265); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20267 = 12'h40b == _T_643 ? $signed(7'shf) : $signed(_GEN_20266); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20268 = 12'h40c == _T_643 ? $signed(7'shf) : $signed(_GEN_20267); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20269 = 12'h40d == _T_643 ? $signed(7'she) : $signed(_GEN_20268); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20270 = 12'h40e == _T_643 ? $signed(7'shd) : $signed(_GEN_20269); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20271 = 12'h40f == _T_643 ? $signed(7'shc) : $signed(_GEN_20270); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20272 = 12'h410 == _T_643 ? $signed(7'shc) : $signed(_GEN_20271); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20273 = 12'h411 == _T_643 ? $signed(7'shb) : $signed(_GEN_20272); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20274 = 12'h412 == _T_643 ? $signed(7'sha) : $signed(_GEN_20273); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20275 = 12'h413 == _T_643 ? $signed(7'sha) : $signed(_GEN_20274); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20276 = 12'h414 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20275); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20277 = 12'h415 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20276); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20278 = 12'h416 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20277); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20279 = 12'h417 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20278); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20280 = 12'h418 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20279); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20281 = 12'h419 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20280); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20282 = 12'h41a == _T_643 ? $signed(7'sh5) : $signed(_GEN_20281); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20283 = 12'h41b == _T_643 ? $signed(7'sh4) : $signed(_GEN_20282); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20284 = 12'h41c == _T_643 ? $signed(7'sh3) : $signed(_GEN_20283); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20285 = 12'h41d == _T_643 ? $signed(7'sh3) : $signed(_GEN_20284); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20286 = 12'h41e == _T_643 ? $signed(7'sh2) : $signed(_GEN_20285); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20287 = 12'h41f == _T_643 ? $signed(7'sh1) : $signed(_GEN_20286); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20288 = 12'h420 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20287); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20289 = 12'h421 == _T_643 ? $signed(7'sh0) : $signed(_GEN_20288); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20290 = 12'h422 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20289); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20291 = 12'h423 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20290); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20292 = 12'h424 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20291); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20293 = 12'h425 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20292); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20294 = 12'h426 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20293); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20295 = 12'h427 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20294); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20296 = 12'h428 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20295); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20297 = 12'h429 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20296); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20298 = 12'h42a == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20297); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20299 = 12'h42b == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20298); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20300 = 12'h42c == _T_643 ? $signed(7'sh19) : $signed(_GEN_20299); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20301 = 12'h42d == _T_643 ? $signed(7'sh18) : $signed(_GEN_20300); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20302 = 12'h42e == _T_643 ? $signed(7'sh18) : $signed(_GEN_20301); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20303 = 12'h42f == _T_643 ? $signed(7'sh17) : $signed(_GEN_20302); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20304 = 12'h430 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20303); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20305 = 12'h431 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20304); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20306 = 12'h432 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20305); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20307 = 12'h433 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20306); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20308 = 12'h434 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20307); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20309 = 12'h435 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20308); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20310 = 12'h436 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20309); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20311 = 12'h437 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20310); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20312 = 12'h438 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20311); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20313 = 12'h439 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20312); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20314 = 12'h43a == _T_643 ? $signed(7'shf) : $signed(_GEN_20313); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20315 = 12'h43b == _T_643 ? $signed(7'shf) : $signed(_GEN_20314); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20316 = 12'h43c == _T_643 ? $signed(7'she) : $signed(_GEN_20315); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20317 = 12'h43d == _T_643 ? $signed(7'shd) : $signed(_GEN_20316); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20318 = 12'h43e == _T_643 ? $signed(7'shc) : $signed(_GEN_20317); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20319 = 12'h43f == _T_643 ? $signed(7'shc) : $signed(_GEN_20318); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20320 = 12'h440 == _T_643 ? $signed(7'shb) : $signed(_GEN_20319); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20321 = 12'h441 == _T_643 ? $signed(7'sha) : $signed(_GEN_20320); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20322 = 12'h442 == _T_643 ? $signed(7'sha) : $signed(_GEN_20321); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20323 = 12'h443 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20322); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20324 = 12'h444 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20323); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20325 = 12'h445 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20324); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20326 = 12'h446 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20325); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20327 = 12'h447 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20326); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20328 = 12'h448 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20327); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20329 = 12'h449 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20328); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20330 = 12'h44a == _T_643 ? $signed(7'sh4) : $signed(_GEN_20329); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20331 = 12'h44b == _T_643 ? $signed(7'sh3) : $signed(_GEN_20330); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20332 = 12'h44c == _T_643 ? $signed(7'sh3) : $signed(_GEN_20331); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20333 = 12'h44d == _T_643 ? $signed(7'sh2) : $signed(_GEN_20332); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20334 = 12'h44e == _T_643 ? $signed(7'sh1) : $signed(_GEN_20333); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20335 = 12'h44f == _T_643 ? $signed(7'sh0) : $signed(_GEN_20334); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20336 = 12'h450 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20335); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20337 = 12'h451 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20336); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20338 = 12'h452 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20337); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20339 = 12'h453 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20338); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20340 = 12'h454 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20339); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20341 = 12'h455 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20340); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20342 = 12'h456 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20341); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20343 = 12'h457 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20342); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20344 = 12'h458 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20343); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20345 = 12'h459 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20344); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20346 = 12'h45a == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20345); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20347 = 12'h45b == _T_643 ? $signed(7'sh19) : $signed(_GEN_20346); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20348 = 12'h45c == _T_643 ? $signed(7'sh18) : $signed(_GEN_20347); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20349 = 12'h45d == _T_643 ? $signed(7'sh18) : $signed(_GEN_20348); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20350 = 12'h45e == _T_643 ? $signed(7'sh17) : $signed(_GEN_20349); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20351 = 12'h45f == _T_643 ? $signed(7'sh16) : $signed(_GEN_20350); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20352 = 12'h460 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20351); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20353 = 12'h461 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20352); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20354 = 12'h462 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20353); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20355 = 12'h463 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20354); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20356 = 12'h464 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20355); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20357 = 12'h465 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20356); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20358 = 12'h466 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20357); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20359 = 12'h467 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20358); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20360 = 12'h468 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20359); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20361 = 12'h469 == _T_643 ? $signed(7'shf) : $signed(_GEN_20360); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20362 = 12'h46a == _T_643 ? $signed(7'shf) : $signed(_GEN_20361); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20363 = 12'h46b == _T_643 ? $signed(7'she) : $signed(_GEN_20362); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20364 = 12'h46c == _T_643 ? $signed(7'shd) : $signed(_GEN_20363); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20365 = 12'h46d == _T_643 ? $signed(7'shc) : $signed(_GEN_20364); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20366 = 12'h46e == _T_643 ? $signed(7'shc) : $signed(_GEN_20365); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20367 = 12'h46f == _T_643 ? $signed(7'shb) : $signed(_GEN_20366); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20368 = 12'h470 == _T_643 ? $signed(7'sha) : $signed(_GEN_20367); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20369 = 12'h471 == _T_643 ? $signed(7'sha) : $signed(_GEN_20368); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20370 = 12'h472 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20369); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20371 = 12'h473 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20370); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20372 = 12'h474 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20371); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20373 = 12'h475 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20372); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20374 = 12'h476 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20373); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20375 = 12'h477 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20374); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20376 = 12'h478 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20375); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20377 = 12'h479 == _T_643 ? $signed(7'sh4) : $signed(_GEN_20376); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20378 = 12'h47a == _T_643 ? $signed(7'sh3) : $signed(_GEN_20377); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20379 = 12'h47b == _T_643 ? $signed(7'sh3) : $signed(_GEN_20378); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20380 = 12'h47c == _T_643 ? $signed(7'sh2) : $signed(_GEN_20379); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20381 = 12'h47d == _T_643 ? $signed(7'sh1) : $signed(_GEN_20380); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20382 = 12'h47e == _T_643 ? $signed(7'sh22) : $signed(_GEN_20381); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20383 = 12'h47f == _T_643 ? $signed(7'sh21) : $signed(_GEN_20382); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20384 = 12'h480 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20383); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20385 = 12'h481 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20384); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20386 = 12'h482 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20385); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20387 = 12'h483 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20386); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20388 = 12'h484 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20387); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20389 = 12'h485 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20388); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20390 = 12'h486 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20389); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20391 = 12'h487 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20390); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20392 = 12'h488 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20391); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20393 = 12'h489 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20392); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20394 = 12'h48a == _T_643 ? $signed(7'sh19) : $signed(_GEN_20393); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20395 = 12'h48b == _T_643 ? $signed(7'sh18) : $signed(_GEN_20394); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20396 = 12'h48c == _T_643 ? $signed(7'sh18) : $signed(_GEN_20395); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20397 = 12'h48d == _T_643 ? $signed(7'sh17) : $signed(_GEN_20396); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20398 = 12'h48e == _T_643 ? $signed(7'sh16) : $signed(_GEN_20397); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20399 = 12'h48f == _T_643 ? $signed(7'sh16) : $signed(_GEN_20398); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20400 = 12'h490 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20399); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20401 = 12'h491 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20400); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20402 = 12'h492 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20401); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20403 = 12'h493 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20402); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20404 = 12'h494 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20403); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20405 = 12'h495 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20404); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20406 = 12'h496 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20405); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20407 = 12'h497 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20406); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20408 = 12'h498 == _T_643 ? $signed(7'shf) : $signed(_GEN_20407); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20409 = 12'h499 == _T_643 ? $signed(7'shf) : $signed(_GEN_20408); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20410 = 12'h49a == _T_643 ? $signed(7'she) : $signed(_GEN_20409); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20411 = 12'h49b == _T_643 ? $signed(7'shd) : $signed(_GEN_20410); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20412 = 12'h49c == _T_643 ? $signed(7'shc) : $signed(_GEN_20411); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20413 = 12'h49d == _T_643 ? $signed(7'shc) : $signed(_GEN_20412); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20414 = 12'h49e == _T_643 ? $signed(7'shb) : $signed(_GEN_20413); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20415 = 12'h49f == _T_643 ? $signed(7'sha) : $signed(_GEN_20414); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20416 = 12'h4a0 == _T_643 ? $signed(7'sha) : $signed(_GEN_20415); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20417 = 12'h4a1 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20416); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20418 = 12'h4a2 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20417); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20419 = 12'h4a3 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20418); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20420 = 12'h4a4 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20419); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20421 = 12'h4a5 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20420); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20422 = 12'h4a6 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20421); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20423 = 12'h4a7 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20422); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20424 = 12'h4a8 == _T_643 ? $signed(7'sh4) : $signed(_GEN_20423); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20425 = 12'h4a9 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20424); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20426 = 12'h4aa == _T_643 ? $signed(7'sh3) : $signed(_GEN_20425); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20427 = 12'h4ab == _T_643 ? $signed(7'sh2) : $signed(_GEN_20426); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20428 = 12'h4ac == _T_643 ? $signed(7'sh22) : $signed(_GEN_20427); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20429 = 12'h4ad == _T_643 ? $signed(7'sh22) : $signed(_GEN_20428); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20430 = 12'h4ae == _T_643 ? $signed(7'sh21) : $signed(_GEN_20429); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20431 = 12'h4af == _T_643 ? $signed(7'sh20) : $signed(_GEN_20430); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20432 = 12'h4b0 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20431); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20433 = 12'h4b1 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20432); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20434 = 12'h4b2 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20433); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20435 = 12'h4b3 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20434); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20436 = 12'h4b4 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20435); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20437 = 12'h4b5 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20436); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20438 = 12'h4b6 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20437); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20439 = 12'h4b7 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20438); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20440 = 12'h4b8 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20439); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20441 = 12'h4b9 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20440); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20442 = 12'h4ba == _T_643 ? $signed(7'sh18) : $signed(_GEN_20441); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20443 = 12'h4bb == _T_643 ? $signed(7'sh18) : $signed(_GEN_20442); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20444 = 12'h4bc == _T_643 ? $signed(7'sh17) : $signed(_GEN_20443); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20445 = 12'h4bd == _T_643 ? $signed(7'sh16) : $signed(_GEN_20444); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20446 = 12'h4be == _T_643 ? $signed(7'sh16) : $signed(_GEN_20445); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20447 = 12'h4bf == _T_643 ? $signed(7'sh15) : $signed(_GEN_20446); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20448 = 12'h4c0 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20447); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20449 = 12'h4c1 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20448); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20450 = 12'h4c2 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20449); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20451 = 12'h4c3 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20450); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20452 = 12'h4c4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20451); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20453 = 12'h4c5 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20452); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20454 = 12'h4c6 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20453); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20455 = 12'h4c7 == _T_643 ? $signed(7'shf) : $signed(_GEN_20454); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20456 = 12'h4c8 == _T_643 ? $signed(7'shf) : $signed(_GEN_20455); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20457 = 12'h4c9 == _T_643 ? $signed(7'she) : $signed(_GEN_20456); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20458 = 12'h4ca == _T_643 ? $signed(7'shd) : $signed(_GEN_20457); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20459 = 12'h4cb == _T_643 ? $signed(7'shc) : $signed(_GEN_20458); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20460 = 12'h4cc == _T_643 ? $signed(7'shc) : $signed(_GEN_20459); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20461 = 12'h4cd == _T_643 ? $signed(7'shb) : $signed(_GEN_20460); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20462 = 12'h4ce == _T_643 ? $signed(7'sha) : $signed(_GEN_20461); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20463 = 12'h4cf == _T_643 ? $signed(7'sha) : $signed(_GEN_20462); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20464 = 12'h4d0 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20463); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20465 = 12'h4d1 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20464); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20466 = 12'h4d2 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20465); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20467 = 12'h4d3 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20466); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20468 = 12'h4d4 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20467); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20469 = 12'h4d5 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20468); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20470 = 12'h4d6 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20469); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20471 = 12'h4d7 == _T_643 ? $signed(7'sh4) : $signed(_GEN_20470); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20472 = 12'h4d8 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20471); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20473 = 12'h4d9 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20472); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20474 = 12'h4da == _T_643 ? $signed(7'sh23) : $signed(_GEN_20473); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20475 = 12'h4db == _T_643 ? $signed(7'sh22) : $signed(_GEN_20474); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20476 = 12'h4dc == _T_643 ? $signed(7'sh22) : $signed(_GEN_20475); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20477 = 12'h4dd == _T_643 ? $signed(7'sh21) : $signed(_GEN_20476); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20478 = 12'h4de == _T_643 ? $signed(7'sh20) : $signed(_GEN_20477); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20479 = 12'h4df == _T_643 ? $signed(7'sh20) : $signed(_GEN_20478); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20480 = 12'h4e0 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20479); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20481 = 12'h4e1 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20480); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20482 = 12'h4e2 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20481); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20483 = 12'h4e3 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20482); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20484 = 12'h4e4 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20483); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20485 = 12'h4e5 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20484); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20486 = 12'h4e6 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20485); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20487 = 12'h4e7 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20486); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20488 = 12'h4e8 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20487); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20489 = 12'h4e9 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20488); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20490 = 12'h4ea == _T_643 ? $signed(7'sh18) : $signed(_GEN_20489); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20491 = 12'h4eb == _T_643 ? $signed(7'sh17) : $signed(_GEN_20490); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20492 = 12'h4ec == _T_643 ? $signed(7'sh16) : $signed(_GEN_20491); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20493 = 12'h4ed == _T_643 ? $signed(7'sh16) : $signed(_GEN_20492); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20494 = 12'h4ee == _T_643 ? $signed(7'sh15) : $signed(_GEN_20493); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20495 = 12'h4ef == _T_643 ? $signed(7'sh14) : $signed(_GEN_20494); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20496 = 12'h4f0 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20495); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20497 = 12'h4f1 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20496); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20498 = 12'h4f2 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20497); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20499 = 12'h4f3 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20498); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20500 = 12'h4f4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20499); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20501 = 12'h4f5 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20500); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20502 = 12'h4f6 == _T_643 ? $signed(7'shf) : $signed(_GEN_20501); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20503 = 12'h4f7 == _T_643 ? $signed(7'shf) : $signed(_GEN_20502); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20504 = 12'h4f8 == _T_643 ? $signed(7'she) : $signed(_GEN_20503); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20505 = 12'h4f9 == _T_643 ? $signed(7'shd) : $signed(_GEN_20504); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20506 = 12'h4fa == _T_643 ? $signed(7'shc) : $signed(_GEN_20505); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20507 = 12'h4fb == _T_643 ? $signed(7'shc) : $signed(_GEN_20506); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20508 = 12'h4fc == _T_643 ? $signed(7'shb) : $signed(_GEN_20507); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20509 = 12'h4fd == _T_643 ? $signed(7'sha) : $signed(_GEN_20508); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20510 = 12'h4fe == _T_643 ? $signed(7'sha) : $signed(_GEN_20509); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20511 = 12'h4ff == _T_643 ? $signed(7'sh9) : $signed(_GEN_20510); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20512 = 12'h500 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20511); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20513 = 12'h501 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20512); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20514 = 12'h502 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20513); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20515 = 12'h503 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20514); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20516 = 12'h504 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20515); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20517 = 12'h505 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20516); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20518 = 12'h506 == _T_643 ? $signed(7'sh4) : $signed(_GEN_20517); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20519 = 12'h507 == _T_643 ? $signed(7'sh3) : $signed(_GEN_20518); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20520 = 12'h508 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20519); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20521 = 12'h509 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20520); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20522 = 12'h50a == _T_643 ? $signed(7'sh22) : $signed(_GEN_20521); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20523 = 12'h50b == _T_643 ? $signed(7'sh22) : $signed(_GEN_20522); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20524 = 12'h50c == _T_643 ? $signed(7'sh21) : $signed(_GEN_20523); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20525 = 12'h50d == _T_643 ? $signed(7'sh20) : $signed(_GEN_20524); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20526 = 12'h50e == _T_643 ? $signed(7'sh20) : $signed(_GEN_20525); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20527 = 12'h50f == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20526); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20528 = 12'h510 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20527); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20529 = 12'h511 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20528); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20530 = 12'h512 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20529); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20531 = 12'h513 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20530); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20532 = 12'h514 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20531); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20533 = 12'h515 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20532); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20534 = 12'h516 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20533); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20535 = 12'h517 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20534); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20536 = 12'h518 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20535); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20537 = 12'h519 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20536); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20538 = 12'h51a == _T_643 ? $signed(7'sh17) : $signed(_GEN_20537); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20539 = 12'h51b == _T_643 ? $signed(7'sh16) : $signed(_GEN_20538); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20540 = 12'h51c == _T_643 ? $signed(7'sh16) : $signed(_GEN_20539); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20541 = 12'h51d == _T_643 ? $signed(7'sh15) : $signed(_GEN_20540); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20542 = 12'h51e == _T_643 ? $signed(7'sh14) : $signed(_GEN_20541); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20543 = 12'h51f == _T_643 ? $signed(7'sh14) : $signed(_GEN_20542); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20544 = 12'h520 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20543); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20545 = 12'h521 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20544); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20546 = 12'h522 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20545); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20547 = 12'h523 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20546); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20548 = 12'h524 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20547); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20549 = 12'h525 == _T_643 ? $signed(7'shf) : $signed(_GEN_20548); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20550 = 12'h526 == _T_643 ? $signed(7'shf) : $signed(_GEN_20549); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20551 = 12'h527 == _T_643 ? $signed(7'she) : $signed(_GEN_20550); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20552 = 12'h528 == _T_643 ? $signed(7'shd) : $signed(_GEN_20551); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20553 = 12'h529 == _T_643 ? $signed(7'shc) : $signed(_GEN_20552); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20554 = 12'h52a == _T_643 ? $signed(7'shc) : $signed(_GEN_20553); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20555 = 12'h52b == _T_643 ? $signed(7'shb) : $signed(_GEN_20554); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20556 = 12'h52c == _T_643 ? $signed(7'sha) : $signed(_GEN_20555); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20557 = 12'h52d == _T_643 ? $signed(7'sha) : $signed(_GEN_20556); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20558 = 12'h52e == _T_643 ? $signed(7'sh9) : $signed(_GEN_20557); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20559 = 12'h52f == _T_643 ? $signed(7'sh8) : $signed(_GEN_20558); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20560 = 12'h530 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20559); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20561 = 12'h531 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20560); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20562 = 12'h532 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20561); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20563 = 12'h533 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20562); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20564 = 12'h534 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20563); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20565 = 12'h535 == _T_643 ? $signed(7'sh4) : $signed(_GEN_20564); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20566 = 12'h536 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20565); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20567 = 12'h537 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20566); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20568 = 12'h538 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20567); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20569 = 12'h539 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20568); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20570 = 12'h53a == _T_643 ? $signed(7'sh22) : $signed(_GEN_20569); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20571 = 12'h53b == _T_643 ? $signed(7'sh21) : $signed(_GEN_20570); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20572 = 12'h53c == _T_643 ? $signed(7'sh20) : $signed(_GEN_20571); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20573 = 12'h53d == _T_643 ? $signed(7'sh20) : $signed(_GEN_20572); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20574 = 12'h53e == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20573); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20575 = 12'h53f == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20574); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20576 = 12'h540 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20575); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20577 = 12'h541 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20576); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20578 = 12'h542 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20577); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20579 = 12'h543 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20578); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20580 = 12'h544 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20579); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20581 = 12'h545 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20580); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20582 = 12'h546 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20581); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20583 = 12'h547 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20582); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20584 = 12'h548 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20583); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20585 = 12'h549 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20584); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20586 = 12'h54a == _T_643 ? $signed(7'sh16) : $signed(_GEN_20585); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20587 = 12'h54b == _T_643 ? $signed(7'sh16) : $signed(_GEN_20586); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20588 = 12'h54c == _T_643 ? $signed(7'sh15) : $signed(_GEN_20587); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20589 = 12'h54d == _T_643 ? $signed(7'sh14) : $signed(_GEN_20588); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20590 = 12'h54e == _T_643 ? $signed(7'sh14) : $signed(_GEN_20589); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20591 = 12'h54f == _T_643 ? $signed(7'sh13) : $signed(_GEN_20590); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20592 = 12'h550 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20591); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20593 = 12'h551 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20592); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20594 = 12'h552 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20593); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20595 = 12'h553 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20594); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20596 = 12'h554 == _T_643 ? $signed(7'shf) : $signed(_GEN_20595); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20597 = 12'h555 == _T_643 ? $signed(7'shf) : $signed(_GEN_20596); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20598 = 12'h556 == _T_643 ? $signed(7'she) : $signed(_GEN_20597); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20599 = 12'h557 == _T_643 ? $signed(7'shd) : $signed(_GEN_20598); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20600 = 12'h558 == _T_643 ? $signed(7'shc) : $signed(_GEN_20599); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20601 = 12'h559 == _T_643 ? $signed(7'shc) : $signed(_GEN_20600); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20602 = 12'h55a == _T_643 ? $signed(7'shb) : $signed(_GEN_20601); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20603 = 12'h55b == _T_643 ? $signed(7'sha) : $signed(_GEN_20602); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20604 = 12'h55c == _T_643 ? $signed(7'sha) : $signed(_GEN_20603); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20605 = 12'h55d == _T_643 ? $signed(7'sh9) : $signed(_GEN_20604); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20606 = 12'h55e == _T_643 ? $signed(7'sh8) : $signed(_GEN_20605); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20607 = 12'h55f == _T_643 ? $signed(7'sh8) : $signed(_GEN_20606); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20608 = 12'h560 == _T_643 ? $signed(7'sh7) : $signed(_GEN_20607); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20609 = 12'h561 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20608); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20610 = 12'h562 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20609); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20611 = 12'h563 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20610); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20612 = 12'h564 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20611); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20613 = 12'h565 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20612); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20614 = 12'h566 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20613); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20615 = 12'h567 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20614); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20616 = 12'h568 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20615); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20617 = 12'h569 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20616); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20618 = 12'h56a == _T_643 ? $signed(7'sh21) : $signed(_GEN_20617); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20619 = 12'h56b == _T_643 ? $signed(7'sh20) : $signed(_GEN_20618); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20620 = 12'h56c == _T_643 ? $signed(7'sh20) : $signed(_GEN_20619); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20621 = 12'h56d == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20620); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20622 = 12'h56e == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20621); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20623 = 12'h56f == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20622); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20624 = 12'h570 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20623); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20625 = 12'h571 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20624); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20626 = 12'h572 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20625); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20627 = 12'h573 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20626); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20628 = 12'h574 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20627); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20629 = 12'h575 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20628); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20630 = 12'h576 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20629); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20631 = 12'h577 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20630); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20632 = 12'h578 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20631); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20633 = 12'h579 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20632); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20634 = 12'h57a == _T_643 ? $signed(7'sh16) : $signed(_GEN_20633); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20635 = 12'h57b == _T_643 ? $signed(7'sh15) : $signed(_GEN_20634); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20636 = 12'h57c == _T_643 ? $signed(7'sh14) : $signed(_GEN_20635); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20637 = 12'h57d == _T_643 ? $signed(7'sh14) : $signed(_GEN_20636); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20638 = 12'h57e == _T_643 ? $signed(7'sh13) : $signed(_GEN_20637); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20639 = 12'h57f == _T_643 ? $signed(7'sh12) : $signed(_GEN_20638); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20640 = 12'h580 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20639); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20641 = 12'h581 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20640); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20642 = 12'h582 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20641); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20643 = 12'h583 == _T_643 ? $signed(7'shf) : $signed(_GEN_20642); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20644 = 12'h584 == _T_643 ? $signed(7'shf) : $signed(_GEN_20643); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20645 = 12'h585 == _T_643 ? $signed(7'she) : $signed(_GEN_20644); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20646 = 12'h586 == _T_643 ? $signed(7'shd) : $signed(_GEN_20645); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20647 = 12'h587 == _T_643 ? $signed(7'shc) : $signed(_GEN_20646); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20648 = 12'h588 == _T_643 ? $signed(7'shc) : $signed(_GEN_20647); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20649 = 12'h589 == _T_643 ? $signed(7'shb) : $signed(_GEN_20648); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20650 = 12'h58a == _T_643 ? $signed(7'sha) : $signed(_GEN_20649); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20651 = 12'h58b == _T_643 ? $signed(7'sha) : $signed(_GEN_20650); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20652 = 12'h58c == _T_643 ? $signed(7'sh9) : $signed(_GEN_20651); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20653 = 12'h58d == _T_643 ? $signed(7'sh8) : $signed(_GEN_20652); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20654 = 12'h58e == _T_643 ? $signed(7'sh8) : $signed(_GEN_20653); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20655 = 12'h58f == _T_643 ? $signed(7'sh7) : $signed(_GEN_20654); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20656 = 12'h590 == _T_643 ? $signed(7'sh6) : $signed(_GEN_20655); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20657 = 12'h591 == _T_643 ? $signed(7'sh5) : $signed(_GEN_20656); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20658 = 12'h592 == _T_643 ? $signed(7'sh26) : $signed(_GEN_20657); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20659 = 12'h593 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20658); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20660 = 12'h594 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20659); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20661 = 12'h595 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20660); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20662 = 12'h596 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20661); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20663 = 12'h597 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20662); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20664 = 12'h598 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20663); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20665 = 12'h599 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20664); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20666 = 12'h59a == _T_643 ? $signed(7'sh20) : $signed(_GEN_20665); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20667 = 12'h59b == _T_643 ? $signed(7'sh20) : $signed(_GEN_20666); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20668 = 12'h59c == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20667); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20669 = 12'h59d == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20668); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20670 = 12'h59e == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20669); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20671 = 12'h59f == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20670); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20672 = 12'h5a0 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20671); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20673 = 12'h5a1 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20672); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20674 = 12'h5a2 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20673); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20675 = 12'h5a3 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20674); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20676 = 12'h5a4 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20675); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20677 = 12'h5a5 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20676); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20678 = 12'h5a6 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20677); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20679 = 12'h5a7 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20678); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20680 = 12'h5a8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20679); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20681 = 12'h5a9 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20680); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20682 = 12'h5aa == _T_643 ? $signed(7'sh15) : $signed(_GEN_20681); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20683 = 12'h5ab == _T_643 ? $signed(7'sh14) : $signed(_GEN_20682); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20684 = 12'h5ac == _T_643 ? $signed(7'sh14) : $signed(_GEN_20683); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20685 = 12'h5ad == _T_643 ? $signed(7'sh13) : $signed(_GEN_20684); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20686 = 12'h5ae == _T_643 ? $signed(7'sh12) : $signed(_GEN_20685); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20687 = 12'h5af == _T_643 ? $signed(7'sh11) : $signed(_GEN_20686); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20688 = 12'h5b0 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20687); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20689 = 12'h5b1 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20688); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20690 = 12'h5b2 == _T_643 ? $signed(7'shf) : $signed(_GEN_20689); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20691 = 12'h5b3 == _T_643 ? $signed(7'shf) : $signed(_GEN_20690); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20692 = 12'h5b4 == _T_643 ? $signed(7'she) : $signed(_GEN_20691); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20693 = 12'h5b5 == _T_643 ? $signed(7'shd) : $signed(_GEN_20692); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20694 = 12'h5b6 == _T_643 ? $signed(7'shc) : $signed(_GEN_20693); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20695 = 12'h5b7 == _T_643 ? $signed(7'shc) : $signed(_GEN_20694); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20696 = 12'h5b8 == _T_643 ? $signed(7'shb) : $signed(_GEN_20695); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20697 = 12'h5b9 == _T_643 ? $signed(7'sha) : $signed(_GEN_20696); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20698 = 12'h5ba == _T_643 ? $signed(7'sha) : $signed(_GEN_20697); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20699 = 12'h5bb == _T_643 ? $signed(7'sh9) : $signed(_GEN_20698); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20700 = 12'h5bc == _T_643 ? $signed(7'sh8) : $signed(_GEN_20699); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20701 = 12'h5bd == _T_643 ? $signed(7'sh8) : $signed(_GEN_20700); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20702 = 12'h5be == _T_643 ? $signed(7'sh7) : $signed(_GEN_20701); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20703 = 12'h5bf == _T_643 ? $signed(7'sh6) : $signed(_GEN_20702); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20704 = 12'h5c0 == _T_643 ? $signed(7'sh27) : $signed(_GEN_20703); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20705 = 12'h5c1 == _T_643 ? $signed(7'sh26) : $signed(_GEN_20704); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20706 = 12'h5c2 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20705); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20707 = 12'h5c3 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20706); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20708 = 12'h5c4 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20707); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20709 = 12'h5c5 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20708); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20710 = 12'h5c6 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20709); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20711 = 12'h5c7 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20710); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20712 = 12'h5c8 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20711); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20713 = 12'h5c9 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20712); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20714 = 12'h5ca == _T_643 ? $signed(7'sh20) : $signed(_GEN_20713); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20715 = 12'h5cb == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20714); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20716 = 12'h5cc == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20715); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20717 = 12'h5cd == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20716); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20718 = 12'h5ce == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20717); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20719 = 12'h5cf == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20718); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20720 = 12'h5d0 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20719); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20721 = 12'h5d1 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20720); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20722 = 12'h5d2 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20721); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20723 = 12'h5d3 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20722); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20724 = 12'h5d4 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20723); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20725 = 12'h5d5 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20724); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20726 = 12'h5d6 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20725); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20727 = 12'h5d7 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20726); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20728 = 12'h5d8 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20727); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20729 = 12'h5d9 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20728); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20730 = 12'h5da == _T_643 ? $signed(7'sh14) : $signed(_GEN_20729); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20731 = 12'h5db == _T_643 ? $signed(7'sh14) : $signed(_GEN_20730); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20732 = 12'h5dc == _T_643 ? $signed(7'sh13) : $signed(_GEN_20731); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20733 = 12'h5dd == _T_643 ? $signed(7'sh12) : $signed(_GEN_20732); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20734 = 12'h5de == _T_643 ? $signed(7'sh11) : $signed(_GEN_20733); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20735 = 12'h5df == _T_643 ? $signed(7'sh11) : $signed(_GEN_20734); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20736 = 12'h5e0 == _T_643 ? $signed(7'sh10) : $signed(_GEN_20735); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20737 = 12'h5e1 == _T_643 ? $signed(7'shf) : $signed(_GEN_20736); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20738 = 12'h5e2 == _T_643 ? $signed(7'shf) : $signed(_GEN_20737); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20739 = 12'h5e3 == _T_643 ? $signed(7'she) : $signed(_GEN_20738); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20740 = 12'h5e4 == _T_643 ? $signed(7'shd) : $signed(_GEN_20739); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20741 = 12'h5e5 == _T_643 ? $signed(7'shc) : $signed(_GEN_20740); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20742 = 12'h5e6 == _T_643 ? $signed(7'shc) : $signed(_GEN_20741); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20743 = 12'h5e7 == _T_643 ? $signed(7'shb) : $signed(_GEN_20742); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20744 = 12'h5e8 == _T_643 ? $signed(7'sha) : $signed(_GEN_20743); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20745 = 12'h5e9 == _T_643 ? $signed(7'sha) : $signed(_GEN_20744); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20746 = 12'h5ea == _T_643 ? $signed(7'sh9) : $signed(_GEN_20745); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20747 = 12'h5eb == _T_643 ? $signed(7'sh8) : $signed(_GEN_20746); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20748 = 12'h5ec == _T_643 ? $signed(7'sh8) : $signed(_GEN_20747); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20749 = 12'h5ed == _T_643 ? $signed(7'sh7) : $signed(_GEN_20748); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20750 = 12'h5ee == _T_643 ? $signed(7'sh27) : $signed(_GEN_20749); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20751 = 12'h5ef == _T_643 ? $signed(7'sh27) : $signed(_GEN_20750); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20752 = 12'h5f0 == _T_643 ? $signed(7'sh26) : $signed(_GEN_20751); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20753 = 12'h5f1 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20752); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20754 = 12'h5f2 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20753); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20755 = 12'h5f3 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20754); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20756 = 12'h5f4 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20755); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20757 = 12'h5f5 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20756); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20758 = 12'h5f6 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20757); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20759 = 12'h5f7 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20758); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20760 = 12'h5f8 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20759); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20761 = 12'h5f9 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20760); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20762 = 12'h5fa == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20761); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20763 = 12'h5fb == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20762); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20764 = 12'h5fc == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20763); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20765 = 12'h5fd == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20764); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20766 = 12'h5fe == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20765); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20767 = 12'h5ff == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20766); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20768 = 12'h600 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20767); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20769 = 12'h601 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20768); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20770 = 12'h602 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20769); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20771 = 12'h603 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20770); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20772 = 12'h604 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20771); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20773 = 12'h605 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20772); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20774 = 12'h606 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20773); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20775 = 12'h607 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20774); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20776 = 12'h608 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20775); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20777 = 12'h609 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20776); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20778 = 12'h60a == _T_643 ? $signed(7'sh14) : $signed(_GEN_20777); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20779 = 12'h60b == _T_643 ? $signed(7'sh13) : $signed(_GEN_20778); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20780 = 12'h60c == _T_643 ? $signed(7'sh12) : $signed(_GEN_20779); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20781 = 12'h60d == _T_643 ? $signed(7'sh11) : $signed(_GEN_20780); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20782 = 12'h60e == _T_643 ? $signed(7'sh11) : $signed(_GEN_20781); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20783 = 12'h60f == _T_643 ? $signed(7'sh10) : $signed(_GEN_20782); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20784 = 12'h610 == _T_643 ? $signed(7'shf) : $signed(_GEN_20783); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20785 = 12'h611 == _T_643 ? $signed(7'shf) : $signed(_GEN_20784); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20786 = 12'h612 == _T_643 ? $signed(7'she) : $signed(_GEN_20785); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20787 = 12'h613 == _T_643 ? $signed(7'shd) : $signed(_GEN_20786); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20788 = 12'h614 == _T_643 ? $signed(7'shc) : $signed(_GEN_20787); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20789 = 12'h615 == _T_643 ? $signed(7'shc) : $signed(_GEN_20788); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20790 = 12'h616 == _T_643 ? $signed(7'shb) : $signed(_GEN_20789); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20791 = 12'h617 == _T_643 ? $signed(7'sha) : $signed(_GEN_20790); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20792 = 12'h618 == _T_643 ? $signed(7'sha) : $signed(_GEN_20791); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20793 = 12'h619 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20792); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20794 = 12'h61a == _T_643 ? $signed(7'sh8) : $signed(_GEN_20793); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20795 = 12'h61b == _T_643 ? $signed(7'sh8) : $signed(_GEN_20794); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20796 = 12'h61c == _T_643 ? $signed(7'sh28) : $signed(_GEN_20795); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20797 = 12'h61d == _T_643 ? $signed(7'sh27) : $signed(_GEN_20796); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20798 = 12'h61e == _T_643 ? $signed(7'sh27) : $signed(_GEN_20797); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20799 = 12'h61f == _T_643 ? $signed(7'sh26) : $signed(_GEN_20798); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20800 = 12'h620 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20799); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20801 = 12'h621 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20800); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20802 = 12'h622 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20801); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20803 = 12'h623 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20802); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20804 = 12'h624 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20803); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20805 = 12'h625 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20804); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20806 = 12'h626 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20805); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20807 = 12'h627 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20806); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20808 = 12'h628 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20807); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20809 = 12'h629 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20808); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20810 = 12'h62a == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20809); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20811 = 12'h62b == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20810); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20812 = 12'h62c == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20811); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20813 = 12'h62d == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20812); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20814 = 12'h62e == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20813); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20815 = 12'h62f == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20814); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20816 = 12'h630 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20815); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20817 = 12'h631 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20816); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20818 = 12'h632 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20817); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20819 = 12'h633 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20818); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20820 = 12'h634 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20819); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20821 = 12'h635 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20820); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20822 = 12'h636 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20821); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20823 = 12'h637 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20822); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20824 = 12'h638 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20823); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20825 = 12'h639 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20824); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20826 = 12'h63a == _T_643 ? $signed(7'sh13) : $signed(_GEN_20825); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20827 = 12'h63b == _T_643 ? $signed(7'sh12) : $signed(_GEN_20826); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20828 = 12'h63c == _T_643 ? $signed(7'sh11) : $signed(_GEN_20827); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20829 = 12'h63d == _T_643 ? $signed(7'sh11) : $signed(_GEN_20828); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20830 = 12'h63e == _T_643 ? $signed(7'sh10) : $signed(_GEN_20829); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20831 = 12'h63f == _T_643 ? $signed(7'shf) : $signed(_GEN_20830); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20832 = 12'h640 == _T_643 ? $signed(7'shf) : $signed(_GEN_20831); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20833 = 12'h641 == _T_643 ? $signed(7'she) : $signed(_GEN_20832); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20834 = 12'h642 == _T_643 ? $signed(7'shd) : $signed(_GEN_20833); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20835 = 12'h643 == _T_643 ? $signed(7'shc) : $signed(_GEN_20834); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20836 = 12'h644 == _T_643 ? $signed(7'shc) : $signed(_GEN_20835); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20837 = 12'h645 == _T_643 ? $signed(7'shb) : $signed(_GEN_20836); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20838 = 12'h646 == _T_643 ? $signed(7'sha) : $signed(_GEN_20837); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20839 = 12'h647 == _T_643 ? $signed(7'sha) : $signed(_GEN_20838); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20840 = 12'h648 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20839); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20841 = 12'h649 == _T_643 ? $signed(7'sh8) : $signed(_GEN_20840); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20842 = 12'h64a == _T_643 ? $signed(7'sh29) : $signed(_GEN_20841); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20843 = 12'h64b == _T_643 ? $signed(7'sh28) : $signed(_GEN_20842); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20844 = 12'h64c == _T_643 ? $signed(7'sh27) : $signed(_GEN_20843); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20845 = 12'h64d == _T_643 ? $signed(7'sh27) : $signed(_GEN_20844); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20846 = 12'h64e == _T_643 ? $signed(7'sh26) : $signed(_GEN_20845); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20847 = 12'h64f == _T_643 ? $signed(7'sh25) : $signed(_GEN_20846); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20848 = 12'h650 == _T_643 ? $signed(7'sh25) : $signed(_GEN_20847); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20849 = 12'h651 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20848); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20850 = 12'h652 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20849); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20851 = 12'h653 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20850); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20852 = 12'h654 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20851); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20853 = 12'h655 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20852); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20854 = 12'h656 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20853); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20855 = 12'h657 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20854); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20856 = 12'h658 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20855); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20857 = 12'h659 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20856); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20858 = 12'h65a == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20857); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20859 = 12'h65b == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20858); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20860 = 12'h65c == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20859); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20861 = 12'h65d == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20860); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20862 = 12'h65e == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20861); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20863 = 12'h65f == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20862); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20864 = 12'h660 == _T_643 ? $signed(7'sh19) : $signed(_GEN_20863); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20865 = 12'h661 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20864); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20866 = 12'h662 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20865); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20867 = 12'h663 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20866); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20868 = 12'h664 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20867); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20869 = 12'h665 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20868); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20870 = 12'h666 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20869); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20871 = 12'h667 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20870); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20872 = 12'h668 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20871); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20873 = 12'h669 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20872); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20874 = 12'h66a == _T_643 ? $signed(7'sh12) : $signed(_GEN_20873); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20875 = 12'h66b == _T_643 ? $signed(7'sh11) : $signed(_GEN_20874); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20876 = 12'h66c == _T_643 ? $signed(7'sh11) : $signed(_GEN_20875); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20877 = 12'h66d == _T_643 ? $signed(7'sh10) : $signed(_GEN_20876); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20878 = 12'h66e == _T_643 ? $signed(7'shf) : $signed(_GEN_20877); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20879 = 12'h66f == _T_643 ? $signed(7'shf) : $signed(_GEN_20878); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20880 = 12'h670 == _T_643 ? $signed(7'she) : $signed(_GEN_20879); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20881 = 12'h671 == _T_643 ? $signed(7'shd) : $signed(_GEN_20880); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20882 = 12'h672 == _T_643 ? $signed(7'shc) : $signed(_GEN_20881); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20883 = 12'h673 == _T_643 ? $signed(7'shc) : $signed(_GEN_20882); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20884 = 12'h674 == _T_643 ? $signed(7'shb) : $signed(_GEN_20883); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20885 = 12'h675 == _T_643 ? $signed(7'sha) : $signed(_GEN_20884); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20886 = 12'h676 == _T_643 ? $signed(7'sha) : $signed(_GEN_20885); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20887 = 12'h677 == _T_643 ? $signed(7'sh9) : $signed(_GEN_20886); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20888 = 12'h678 == _T_643 ? $signed(7'sh29) : $signed(_GEN_20887); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20889 = 12'h679 == _T_643 ? $signed(7'sh29) : $signed(_GEN_20888); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20890 = 12'h67a == _T_643 ? $signed(7'sh28) : $signed(_GEN_20889); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20891 = 12'h67b == _T_643 ? $signed(7'sh27) : $signed(_GEN_20890); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20892 = 12'h67c == _T_643 ? $signed(7'sh27) : $signed(_GEN_20891); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20893 = 12'h67d == _T_643 ? $signed(7'sh26) : $signed(_GEN_20892); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20894 = 12'h67e == _T_643 ? $signed(7'sh25) : $signed(_GEN_20893); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20895 = 12'h67f == _T_643 ? $signed(7'sh25) : $signed(_GEN_20894); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20896 = 12'h680 == _T_643 ? $signed(7'sh24) : $signed(_GEN_20895); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20897 = 12'h681 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20896); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20898 = 12'h682 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20897); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20899 = 12'h683 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20898); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20900 = 12'h684 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20899); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20901 = 12'h685 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20900); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20902 = 12'h686 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20901); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20903 = 12'h687 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20902); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20904 = 12'h688 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20903); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20905 = 12'h689 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20904); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20906 = 12'h68a == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20905); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20907 = 12'h68b == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20906); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20908 = 12'h68c == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20907); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20909 = 12'h68d == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20908); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20910 = 12'h68e == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20909); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20911 = 12'h68f == _T_643 ? $signed(7'sh19) : $signed(_GEN_20910); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20912 = 12'h690 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20911); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20913 = 12'h691 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20912); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20914 = 12'h692 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20913); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20915 = 12'h693 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20914); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20916 = 12'h694 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20915); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20917 = 12'h695 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20916); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20918 = 12'h696 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20917); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20919 = 12'h697 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20918); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20920 = 12'h698 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20919); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20921 = 12'h699 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20920); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20922 = 12'h69a == _T_643 ? $signed(7'sh11) : $signed(_GEN_20921); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20923 = 12'h69b == _T_643 ? $signed(7'sh11) : $signed(_GEN_20922); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20924 = 12'h69c == _T_643 ? $signed(7'sh10) : $signed(_GEN_20923); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20925 = 12'h69d == _T_643 ? $signed(7'shf) : $signed(_GEN_20924); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20926 = 12'h69e == _T_643 ? $signed(7'shf) : $signed(_GEN_20925); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20927 = 12'h69f == _T_643 ? $signed(7'she) : $signed(_GEN_20926); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20928 = 12'h6a0 == _T_643 ? $signed(7'shd) : $signed(_GEN_20927); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20929 = 12'h6a1 == _T_643 ? $signed(7'shc) : $signed(_GEN_20928); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20930 = 12'h6a2 == _T_643 ? $signed(7'shc) : $signed(_GEN_20929); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20931 = 12'h6a3 == _T_643 ? $signed(7'shb) : $signed(_GEN_20930); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20932 = 12'h6a4 == _T_643 ? $signed(7'sha) : $signed(_GEN_20931); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20933 = 12'h6a5 == _T_643 ? $signed(7'sha) : $signed(_GEN_20932); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20934 = 12'h6a6 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_20933); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20935 = 12'h6a7 == _T_643 ? $signed(7'sh29) : $signed(_GEN_20934); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20936 = 12'h6a8 == _T_643 ? $signed(7'sh29) : $signed(_GEN_20935); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20937 = 12'h6a9 == _T_643 ? $signed(7'sh28) : $signed(_GEN_20936); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20938 = 12'h6aa == _T_643 ? $signed(7'sh27) : $signed(_GEN_20937); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20939 = 12'h6ab == _T_643 ? $signed(7'sh27) : $signed(_GEN_20938); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20940 = 12'h6ac == _T_643 ? $signed(7'sh26) : $signed(_GEN_20939); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20941 = 12'h6ad == _T_643 ? $signed(7'sh25) : $signed(_GEN_20940); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20942 = 12'h6ae == _T_643 ? $signed(7'sh25) : $signed(_GEN_20941); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20943 = 12'h6af == _T_643 ? $signed(7'sh24) : $signed(_GEN_20942); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20944 = 12'h6b0 == _T_643 ? $signed(7'sh23) : $signed(_GEN_20943); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20945 = 12'h6b1 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20944); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20946 = 12'h6b2 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20945); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20947 = 12'h6b3 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20946); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20948 = 12'h6b4 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20947); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20949 = 12'h6b5 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20948); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20950 = 12'h6b6 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20949); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20951 = 12'h6b7 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20950); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20952 = 12'h6b8 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20951); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20953 = 12'h6b9 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20952); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20954 = 12'h6ba == _T_643 ? $signed(7'sh1c) : $signed(_GEN_20953); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20955 = 12'h6bb == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20954); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20956 = 12'h6bc == _T_643 ? $signed(7'sh1b) : $signed(_GEN_20955); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20957 = 12'h6bd == _T_643 ? $signed(7'sh1a) : $signed(_GEN_20956); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20958 = 12'h6be == _T_643 ? $signed(7'sh19) : $signed(_GEN_20957); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20959 = 12'h6bf == _T_643 ? $signed(7'sh18) : $signed(_GEN_20958); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20960 = 12'h6c0 == _T_643 ? $signed(7'sh18) : $signed(_GEN_20959); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20961 = 12'h6c1 == _T_643 ? $signed(7'sh17) : $signed(_GEN_20960); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20962 = 12'h6c2 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20961); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20963 = 12'h6c3 == _T_643 ? $signed(7'sh16) : $signed(_GEN_20962); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20964 = 12'h6c4 == _T_643 ? $signed(7'sh15) : $signed(_GEN_20963); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20965 = 12'h6c5 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20964); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20966 = 12'h6c6 == _T_643 ? $signed(7'sh14) : $signed(_GEN_20965); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20967 = 12'h6c7 == _T_643 ? $signed(7'sh13) : $signed(_GEN_20966); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20968 = 12'h6c8 == _T_643 ? $signed(7'sh12) : $signed(_GEN_20967); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20969 = 12'h6c9 == _T_643 ? $signed(7'sh11) : $signed(_GEN_20968); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20970 = 12'h6ca == _T_643 ? $signed(7'sh11) : $signed(_GEN_20969); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20971 = 12'h6cb == _T_643 ? $signed(7'sh10) : $signed(_GEN_20970); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20972 = 12'h6cc == _T_643 ? $signed(7'shf) : $signed(_GEN_20971); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20973 = 12'h6cd == _T_643 ? $signed(7'shf) : $signed(_GEN_20972); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20974 = 12'h6ce == _T_643 ? $signed(7'she) : $signed(_GEN_20973); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20975 = 12'h6cf == _T_643 ? $signed(7'shd) : $signed(_GEN_20974); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20976 = 12'h6d0 == _T_643 ? $signed(7'shc) : $signed(_GEN_20975); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20977 = 12'h6d1 == _T_643 ? $signed(7'shc) : $signed(_GEN_20976); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20978 = 12'h6d2 == _T_643 ? $signed(7'shb) : $signed(_GEN_20977); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20979 = 12'h6d3 == _T_643 ? $signed(7'sha) : $signed(_GEN_20978); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20980 = 12'h6d4 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_20979); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20981 = 12'h6d5 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_20980); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20982 = 12'h6d6 == _T_643 ? $signed(7'sh29) : $signed(_GEN_20981); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20983 = 12'h6d7 == _T_643 ? $signed(7'sh29) : $signed(_GEN_20982); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20984 = 12'h6d8 == _T_643 ? $signed(7'sh28) : $signed(_GEN_20983); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20985 = 12'h6d9 == _T_643 ? $signed(7'sh27) : $signed(_GEN_20984); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20986 = 12'h6da == _T_643 ? $signed(7'sh27) : $signed(_GEN_20985); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20987 = 12'h6db == _T_643 ? $signed(7'sh26) : $signed(_GEN_20986); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20988 = 12'h6dc == _T_643 ? $signed(7'sh25) : $signed(_GEN_20987); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20989 = 12'h6dd == _T_643 ? $signed(7'sh25) : $signed(_GEN_20988); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20990 = 12'h6de == _T_643 ? $signed(7'sh24) : $signed(_GEN_20989); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20991 = 12'h6df == _T_643 ? $signed(7'sh23) : $signed(_GEN_20990); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20992 = 12'h6e0 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20991); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20993 = 12'h6e1 == _T_643 ? $signed(7'sh22) : $signed(_GEN_20992); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20994 = 12'h6e2 == _T_643 ? $signed(7'sh21) : $signed(_GEN_20993); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20995 = 12'h6e3 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20994); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20996 = 12'h6e4 == _T_643 ? $signed(7'sh20) : $signed(_GEN_20995); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20997 = 12'h6e5 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_20996); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20998 = 12'h6e6 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_20997); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_20999 = 12'h6e7 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20998); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21000 = 12'h6e8 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_20999); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21001 = 12'h6e9 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21000); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21002 = 12'h6ea == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21001); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21003 = 12'h6eb == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21002); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21004 = 12'h6ec == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21003); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21005 = 12'h6ed == _T_643 ? $signed(7'sh19) : $signed(_GEN_21004); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21006 = 12'h6ee == _T_643 ? $signed(7'sh18) : $signed(_GEN_21005); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21007 = 12'h6ef == _T_643 ? $signed(7'sh18) : $signed(_GEN_21006); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21008 = 12'h6f0 == _T_643 ? $signed(7'sh17) : $signed(_GEN_21007); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21009 = 12'h6f1 == _T_643 ? $signed(7'sh16) : $signed(_GEN_21008); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21010 = 12'h6f2 == _T_643 ? $signed(7'sh16) : $signed(_GEN_21009); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21011 = 12'h6f3 == _T_643 ? $signed(7'sh15) : $signed(_GEN_21010); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21012 = 12'h6f4 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21011); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21013 = 12'h6f5 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21012); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21014 = 12'h6f6 == _T_643 ? $signed(7'sh13) : $signed(_GEN_21013); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21015 = 12'h6f7 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21014); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21016 = 12'h6f8 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21015); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21017 = 12'h6f9 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21016); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21018 = 12'h6fa == _T_643 ? $signed(7'sh10) : $signed(_GEN_21017); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21019 = 12'h6fb == _T_643 ? $signed(7'shf) : $signed(_GEN_21018); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21020 = 12'h6fc == _T_643 ? $signed(7'shf) : $signed(_GEN_21019); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21021 = 12'h6fd == _T_643 ? $signed(7'she) : $signed(_GEN_21020); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21022 = 12'h6fe == _T_643 ? $signed(7'shd) : $signed(_GEN_21021); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21023 = 12'h6ff == _T_643 ? $signed(7'shc) : $signed(_GEN_21022); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21024 = 12'h700 == _T_643 ? $signed(7'shc) : $signed(_GEN_21023); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21025 = 12'h701 == _T_643 ? $signed(7'shb) : $signed(_GEN_21024); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21026 = 12'h702 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21025); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21027 = 12'h703 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_21026); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21028 = 12'h704 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_21027); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21029 = 12'h705 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21028); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21030 = 12'h706 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21029); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21031 = 12'h707 == _T_643 ? $signed(7'sh28) : $signed(_GEN_21030); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21032 = 12'h708 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21031); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21033 = 12'h709 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21032); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21034 = 12'h70a == _T_643 ? $signed(7'sh26) : $signed(_GEN_21033); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21035 = 12'h70b == _T_643 ? $signed(7'sh25) : $signed(_GEN_21034); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21036 = 12'h70c == _T_643 ? $signed(7'sh25) : $signed(_GEN_21035); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21037 = 12'h70d == _T_643 ? $signed(7'sh24) : $signed(_GEN_21036); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21038 = 12'h70e == _T_643 ? $signed(7'sh23) : $signed(_GEN_21037); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21039 = 12'h70f == _T_643 ? $signed(7'sh22) : $signed(_GEN_21038); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21040 = 12'h710 == _T_643 ? $signed(7'sh22) : $signed(_GEN_21039); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21041 = 12'h711 == _T_643 ? $signed(7'sh21) : $signed(_GEN_21040); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21042 = 12'h712 == _T_643 ? $signed(7'sh20) : $signed(_GEN_21041); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21043 = 12'h713 == _T_643 ? $signed(7'sh20) : $signed(_GEN_21042); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21044 = 12'h714 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_21043); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21045 = 12'h715 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_21044); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21046 = 12'h716 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21045); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21047 = 12'h717 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21046); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21048 = 12'h718 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21047); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21049 = 12'h719 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21048); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21050 = 12'h71a == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21049); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21051 = 12'h71b == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21050); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21052 = 12'h71c == _T_643 ? $signed(7'sh19) : $signed(_GEN_21051); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21053 = 12'h71d == _T_643 ? $signed(7'sh18) : $signed(_GEN_21052); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21054 = 12'h71e == _T_643 ? $signed(7'sh18) : $signed(_GEN_21053); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21055 = 12'h71f == _T_643 ? $signed(7'sh17) : $signed(_GEN_21054); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21056 = 12'h720 == _T_643 ? $signed(7'sh16) : $signed(_GEN_21055); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21057 = 12'h721 == _T_643 ? $signed(7'sh16) : $signed(_GEN_21056); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21058 = 12'h722 == _T_643 ? $signed(7'sh15) : $signed(_GEN_21057); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21059 = 12'h723 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21058); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21060 = 12'h724 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21059); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21061 = 12'h725 == _T_643 ? $signed(7'sh13) : $signed(_GEN_21060); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21062 = 12'h726 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21061); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21063 = 12'h727 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21062); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21064 = 12'h728 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21063); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21065 = 12'h729 == _T_643 ? $signed(7'sh10) : $signed(_GEN_21064); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21066 = 12'h72a == _T_643 ? $signed(7'shf) : $signed(_GEN_21065); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21067 = 12'h72b == _T_643 ? $signed(7'shf) : $signed(_GEN_21066); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21068 = 12'h72c == _T_643 ? $signed(7'she) : $signed(_GEN_21067); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21069 = 12'h72d == _T_643 ? $signed(7'shd) : $signed(_GEN_21068); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21070 = 12'h72e == _T_643 ? $signed(7'shc) : $signed(_GEN_21069); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21071 = 12'h72f == _T_643 ? $signed(7'shc) : $signed(_GEN_21070); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21072 = 12'h730 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21071); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21073 = 12'h731 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21072); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21074 = 12'h732 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_21073); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21075 = 12'h733 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_21074); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21076 = 12'h734 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21075); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21077 = 12'h735 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21076); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21078 = 12'h736 == _T_643 ? $signed(7'sh28) : $signed(_GEN_21077); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21079 = 12'h737 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21078); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21080 = 12'h738 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21079); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21081 = 12'h739 == _T_643 ? $signed(7'sh26) : $signed(_GEN_21080); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21082 = 12'h73a == _T_643 ? $signed(7'sh25) : $signed(_GEN_21081); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21083 = 12'h73b == _T_643 ? $signed(7'sh25) : $signed(_GEN_21082); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21084 = 12'h73c == _T_643 ? $signed(7'sh24) : $signed(_GEN_21083); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21085 = 12'h73d == _T_643 ? $signed(7'sh23) : $signed(_GEN_21084); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21086 = 12'h73e == _T_643 ? $signed(7'sh22) : $signed(_GEN_21085); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21087 = 12'h73f == _T_643 ? $signed(7'sh22) : $signed(_GEN_21086); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21088 = 12'h740 == _T_643 ? $signed(7'sh21) : $signed(_GEN_21087); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21089 = 12'h741 == _T_643 ? $signed(7'sh20) : $signed(_GEN_21088); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21090 = 12'h742 == _T_643 ? $signed(7'sh20) : $signed(_GEN_21089); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21091 = 12'h743 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_21090); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21092 = 12'h744 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_21091); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21093 = 12'h745 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21092); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21094 = 12'h746 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21093); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21095 = 12'h747 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21094); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21096 = 12'h748 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21095); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21097 = 12'h749 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21096); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21098 = 12'h74a == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21097); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21099 = 12'h74b == _T_643 ? $signed(7'sh19) : $signed(_GEN_21098); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21100 = 12'h74c == _T_643 ? $signed(7'sh18) : $signed(_GEN_21099); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21101 = 12'h74d == _T_643 ? $signed(7'sh18) : $signed(_GEN_21100); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21102 = 12'h74e == _T_643 ? $signed(7'sh17) : $signed(_GEN_21101); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21103 = 12'h74f == _T_643 ? $signed(7'sh16) : $signed(_GEN_21102); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21104 = 12'h750 == _T_643 ? $signed(7'sh16) : $signed(_GEN_21103); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21105 = 12'h751 == _T_643 ? $signed(7'sh15) : $signed(_GEN_21104); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21106 = 12'h752 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21105); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21107 = 12'h753 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21106); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21108 = 12'h754 == _T_643 ? $signed(7'sh13) : $signed(_GEN_21107); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21109 = 12'h755 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21108); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21110 = 12'h756 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21109); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21111 = 12'h757 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21110); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21112 = 12'h758 == _T_643 ? $signed(7'sh10) : $signed(_GEN_21111); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21113 = 12'h759 == _T_643 ? $signed(7'shf) : $signed(_GEN_21112); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21114 = 12'h75a == _T_643 ? $signed(7'shf) : $signed(_GEN_21113); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21115 = 12'h75b == _T_643 ? $signed(7'she) : $signed(_GEN_21114); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21116 = 12'h75c == _T_643 ? $signed(7'shd) : $signed(_GEN_21115); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21117 = 12'h75d == _T_643 ? $signed(7'shc) : $signed(_GEN_21116); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21118 = 12'h75e == _T_643 ? $signed(7'sh2d) : $signed(_GEN_21117); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21119 = 12'h75f == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21118); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21120 = 12'h760 == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21119); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21121 = 12'h761 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_21120); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21122 = 12'h762 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_21121); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21123 = 12'h763 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21122); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21124 = 12'h764 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21123); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21125 = 12'h765 == _T_643 ? $signed(7'sh28) : $signed(_GEN_21124); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21126 = 12'h766 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21125); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21127 = 12'h767 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21126); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21128 = 12'h768 == _T_643 ? $signed(7'sh26) : $signed(_GEN_21127); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21129 = 12'h769 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21128); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21130 = 12'h76a == _T_643 ? $signed(7'sh25) : $signed(_GEN_21129); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21131 = 12'h76b == _T_643 ? $signed(7'sh24) : $signed(_GEN_21130); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21132 = 12'h76c == _T_643 ? $signed(7'sh23) : $signed(_GEN_21131); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21133 = 12'h76d == _T_643 ? $signed(7'sh22) : $signed(_GEN_21132); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21134 = 12'h76e == _T_643 ? $signed(7'sh22) : $signed(_GEN_21133); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21135 = 12'h76f == _T_643 ? $signed(7'sh21) : $signed(_GEN_21134); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21136 = 12'h770 == _T_643 ? $signed(7'sh20) : $signed(_GEN_21135); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21137 = 12'h771 == _T_643 ? $signed(7'sh20) : $signed(_GEN_21136); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21138 = 12'h772 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_21137); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21139 = 12'h773 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_21138); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21140 = 12'h774 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21139); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21141 = 12'h775 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21140); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21142 = 12'h776 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21141); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21143 = 12'h777 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21142); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21144 = 12'h778 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21143); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21145 = 12'h779 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21144); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21146 = 12'h77a == _T_643 ? $signed(7'sh19) : $signed(_GEN_21145); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21147 = 12'h77b == _T_643 ? $signed(7'sh18) : $signed(_GEN_21146); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21148 = 12'h77c == _T_643 ? $signed(7'sh18) : $signed(_GEN_21147); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21149 = 12'h77d == _T_643 ? $signed(7'sh17) : $signed(_GEN_21148); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21150 = 12'h77e == _T_643 ? $signed(7'sh16) : $signed(_GEN_21149); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21151 = 12'h77f == _T_643 ? $signed(7'sh16) : $signed(_GEN_21150); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21152 = 12'h780 == _T_643 ? $signed(7'sh15) : $signed(_GEN_21151); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21153 = 12'h781 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21152); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21154 = 12'h782 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21153); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21155 = 12'h783 == _T_643 ? $signed(7'sh13) : $signed(_GEN_21154); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21156 = 12'h784 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21155); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21157 = 12'h785 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21156); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21158 = 12'h786 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21157); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21159 = 12'h787 == _T_643 ? $signed(7'sh10) : $signed(_GEN_21158); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21160 = 12'h788 == _T_643 ? $signed(7'shf) : $signed(_GEN_21159); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21161 = 12'h789 == _T_643 ? $signed(7'shf) : $signed(_GEN_21160); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21162 = 12'h78a == _T_643 ? $signed(7'she) : $signed(_GEN_21161); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21163 = 12'h78b == _T_643 ? $signed(7'shd) : $signed(_GEN_21162); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21164 = 12'h78c == _T_643 ? $signed(7'sh2e) : $signed(_GEN_21163); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21165 = 12'h78d == _T_643 ? $signed(7'sh2d) : $signed(_GEN_21164); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21166 = 12'h78e == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21165); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21167 = 12'h78f == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21166); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21168 = 12'h790 == _T_643 ? $signed(7'sh2b) : $signed(_GEN_21167); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21169 = 12'h791 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_21168); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21170 = 12'h792 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21169); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21171 = 12'h793 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21170); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21172 = 12'h794 == _T_643 ? $signed(7'sh28) : $signed(_GEN_21171); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21173 = 12'h795 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21172); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21174 = 12'h796 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21173); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21175 = 12'h797 == _T_643 ? $signed(7'sh26) : $signed(_GEN_21174); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21176 = 12'h798 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21175); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21177 = 12'h799 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21176); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21178 = 12'h79a == _T_643 ? $signed(7'sh24) : $signed(_GEN_21177); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21179 = 12'h79b == _T_643 ? $signed(7'sh23) : $signed(_GEN_21178); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21180 = 12'h79c == _T_643 ? $signed(7'sh22) : $signed(_GEN_21179); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21181 = 12'h79d == _T_643 ? $signed(7'sh22) : $signed(_GEN_21180); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21182 = 12'h79e == _T_643 ? $signed(7'sh21) : $signed(_GEN_21181); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21183 = 12'h79f == _T_643 ? $signed(7'sh20) : $signed(_GEN_21182); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21184 = 12'h7a0 == _T_643 ? $signed(7'sh20) : $signed(_GEN_21183); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21185 = 12'h7a1 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_21184); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21186 = 12'h7a2 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_21185); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21187 = 12'h7a3 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21186); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21188 = 12'h7a4 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21187); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21189 = 12'h7a5 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21188); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21190 = 12'h7a6 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21189); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21191 = 12'h7a7 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21190); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21192 = 12'h7a8 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21191); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21193 = 12'h7a9 == _T_643 ? $signed(7'sh19) : $signed(_GEN_21192); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21194 = 12'h7aa == _T_643 ? $signed(7'sh18) : $signed(_GEN_21193); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21195 = 12'h7ab == _T_643 ? $signed(7'sh18) : $signed(_GEN_21194); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21196 = 12'h7ac == _T_643 ? $signed(7'sh17) : $signed(_GEN_21195); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21197 = 12'h7ad == _T_643 ? $signed(7'sh16) : $signed(_GEN_21196); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21198 = 12'h7ae == _T_643 ? $signed(7'sh16) : $signed(_GEN_21197); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21199 = 12'h7af == _T_643 ? $signed(7'sh15) : $signed(_GEN_21198); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21200 = 12'h7b0 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21199); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21201 = 12'h7b1 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21200); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21202 = 12'h7b2 == _T_643 ? $signed(7'sh13) : $signed(_GEN_21201); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21203 = 12'h7b3 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21202); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21204 = 12'h7b4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21203); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21205 = 12'h7b5 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21204); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21206 = 12'h7b6 == _T_643 ? $signed(7'sh10) : $signed(_GEN_21205); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21207 = 12'h7b7 == _T_643 ? $signed(7'shf) : $signed(_GEN_21206); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21208 = 12'h7b8 == _T_643 ? $signed(7'shf) : $signed(_GEN_21207); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21209 = 12'h7b9 == _T_643 ? $signed(7'she) : $signed(_GEN_21208); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21210 = 12'h7ba == _T_643 ? $signed(7'sh2e) : $signed(_GEN_21209); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21211 = 12'h7bb == _T_643 ? $signed(7'sh2e) : $signed(_GEN_21210); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21212 = 12'h7bc == _T_643 ? $signed(7'sh2d) : $signed(_GEN_21211); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21213 = 12'h7bd == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21212); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21214 = 12'h7be == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21213); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21215 = 12'h7bf == _T_643 ? $signed(7'sh2b) : $signed(_GEN_21214); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21216 = 12'h7c0 == _T_643 ? $signed(7'sh2a) : $signed(_GEN_21215); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21217 = 12'h7c1 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21216); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21218 = 12'h7c2 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21217); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21219 = 12'h7c3 == _T_643 ? $signed(7'sh28) : $signed(_GEN_21218); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21220 = 12'h7c4 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21219); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21221 = 12'h7c5 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21220); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21222 = 12'h7c6 == _T_643 ? $signed(7'sh26) : $signed(_GEN_21221); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21223 = 12'h7c7 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21222); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21224 = 12'h7c8 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21223); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21225 = 12'h7c9 == _T_643 ? $signed(7'sh24) : $signed(_GEN_21224); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21226 = 12'h7ca == _T_643 ? $signed(7'sh23) : $signed(_GEN_21225); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21227 = 12'h7cb == _T_643 ? $signed(7'sh22) : $signed(_GEN_21226); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21228 = 12'h7cc == _T_643 ? $signed(7'sh22) : $signed(_GEN_21227); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21229 = 12'h7cd == _T_643 ? $signed(7'sh21) : $signed(_GEN_21228); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21230 = 12'h7ce == _T_643 ? $signed(7'sh20) : $signed(_GEN_21229); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21231 = 12'h7cf == _T_643 ? $signed(7'sh20) : $signed(_GEN_21230); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21232 = 12'h7d0 == _T_643 ? $signed(7'sh1f) : $signed(_GEN_21231); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21233 = 12'h7d1 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_21232); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21234 = 12'h7d2 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21233); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21235 = 12'h7d3 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21234); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21236 = 12'h7d4 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21235); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21237 = 12'h7d5 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21236); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21238 = 12'h7d6 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21237); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21239 = 12'h7d7 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21238); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21240 = 12'h7d8 == _T_643 ? $signed(7'sh19) : $signed(_GEN_21239); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21241 = 12'h7d9 == _T_643 ? $signed(7'sh18) : $signed(_GEN_21240); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21242 = 12'h7da == _T_643 ? $signed(7'sh18) : $signed(_GEN_21241); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21243 = 12'h7db == _T_643 ? $signed(7'sh17) : $signed(_GEN_21242); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21244 = 12'h7dc == _T_643 ? $signed(7'sh16) : $signed(_GEN_21243); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21245 = 12'h7dd == _T_643 ? $signed(7'sh16) : $signed(_GEN_21244); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21246 = 12'h7de == _T_643 ? $signed(7'sh15) : $signed(_GEN_21245); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21247 = 12'h7df == _T_643 ? $signed(7'sh14) : $signed(_GEN_21246); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21248 = 12'h7e0 == _T_643 ? $signed(7'sh14) : $signed(_GEN_21247); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21249 = 12'h7e1 == _T_643 ? $signed(7'sh13) : $signed(_GEN_21248); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21250 = 12'h7e2 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21249); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21251 = 12'h7e3 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21250); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21252 = 12'h7e4 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21251); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21253 = 12'h7e5 == _T_643 ? $signed(7'sh10) : $signed(_GEN_21252); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21254 = 12'h7e6 == _T_643 ? $signed(7'shf) : $signed(_GEN_21253); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21255 = 12'h7e7 == _T_643 ? $signed(7'shf) : $signed(_GEN_21254); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21256 = 12'h7e8 == _T_643 ? $signed(7'sh2f) : $signed(_GEN_21255); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21257 = 12'h7e9 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_21256); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21258 = 12'h7ea == _T_643 ? $signed(7'sh2e) : $signed(_GEN_21257); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21259 = 12'h7eb == _T_643 ? $signed(7'sh2d) : $signed(_GEN_21258); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21260 = 12'h7ec == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21259); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21261 = 12'h7ed == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21260); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21262 = 12'h7ee == _T_643 ? $signed(7'sh2b) : $signed(_GEN_21261); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21263 = 12'h7ef == _T_643 ? $signed(7'sh2a) : $signed(_GEN_21262); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21264 = 12'h7f0 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21263); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21265 = 12'h7f1 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21264); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21266 = 12'h7f2 == _T_643 ? $signed(7'sh28) : $signed(_GEN_21265); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21267 = 12'h7f3 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21266); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21268 = 12'h7f4 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21267); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21269 = 12'h7f5 == _T_643 ? $signed(7'sh26) : $signed(_GEN_21268); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21270 = 12'h7f6 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21269); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21271 = 12'h7f7 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21270); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21272 = 12'h7f8 == _T_643 ? $signed(7'sh24) : $signed(_GEN_21271); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21273 = 12'h7f9 == _T_643 ? $signed(7'sh23) : $signed(_GEN_21272); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21274 = 12'h7fa == _T_643 ? $signed(7'sh22) : $signed(_GEN_21273); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21275 = 12'h7fb == _T_643 ? $signed(7'sh22) : $signed(_GEN_21274); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21276 = 12'h7fc == _T_643 ? $signed(7'sh21) : $signed(_GEN_21275); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21277 = 12'h7fd == _T_643 ? $signed(7'sh20) : $signed(_GEN_21276); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21278 = 12'h7fe == _T_643 ? $signed(7'sh20) : $signed(_GEN_21277); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21279 = 12'h7ff == _T_643 ? $signed(7'sh1f) : $signed(_GEN_21278); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21280 = 12'h800 == _T_643 ? $signed(7'sh1e) : $signed(_GEN_21279); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21281 = 12'h801 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21280); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21282 = 12'h802 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21281); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21283 = 12'h803 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21282); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21284 = 12'h804 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21283); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21285 = 12'h805 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21284); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21286 = 12'h806 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21285); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21287 = 12'h807 == _T_643 ? $signed(7'sh19) : $signed(_GEN_21286); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21288 = 12'h808 == _T_643 ? $signed(7'sh18) : $signed(_GEN_21287); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21289 = 12'h809 == _T_643 ? $signed(7'sh18) : $signed(_GEN_21288); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21290 = 12'h80a == _T_643 ? $signed(7'sh17) : $signed(_GEN_21289); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21291 = 12'h80b == _T_643 ? $signed(7'sh16) : $signed(_GEN_21290); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21292 = 12'h80c == _T_643 ? $signed(7'sh16) : $signed(_GEN_21291); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21293 = 12'h80d == _T_643 ? $signed(7'sh15) : $signed(_GEN_21292); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21294 = 12'h80e == _T_643 ? $signed(7'sh14) : $signed(_GEN_21293); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21295 = 12'h80f == _T_643 ? $signed(7'sh14) : $signed(_GEN_21294); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21296 = 12'h810 == _T_643 ? $signed(7'sh13) : $signed(_GEN_21295); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21297 = 12'h811 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21296); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21298 = 12'h812 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21297); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21299 = 12'h813 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21298); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21300 = 12'h814 == _T_643 ? $signed(7'sh10) : $signed(_GEN_21299); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21301 = 12'h815 == _T_643 ? $signed(7'shf) : $signed(_GEN_21300); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21302 = 12'h816 == _T_643 ? $signed(7'sh30) : $signed(_GEN_21301); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21303 = 12'h817 == _T_643 ? $signed(7'sh2f) : $signed(_GEN_21302); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21304 = 12'h818 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_21303); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21305 = 12'h819 == _T_643 ? $signed(7'sh2e) : $signed(_GEN_21304); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21306 = 12'h81a == _T_643 ? $signed(7'sh2d) : $signed(_GEN_21305); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21307 = 12'h81b == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21306); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21308 = 12'h81c == _T_643 ? $signed(7'sh2c) : $signed(_GEN_21307); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21309 = 12'h81d == _T_643 ? $signed(7'sh2b) : $signed(_GEN_21308); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21310 = 12'h81e == _T_643 ? $signed(7'sh2a) : $signed(_GEN_21309); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21311 = 12'h81f == _T_643 ? $signed(7'sh29) : $signed(_GEN_21310); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21312 = 12'h820 == _T_643 ? $signed(7'sh29) : $signed(_GEN_21311); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21313 = 12'h821 == _T_643 ? $signed(7'sh28) : $signed(_GEN_21312); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21314 = 12'h822 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21313); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21315 = 12'h823 == _T_643 ? $signed(7'sh27) : $signed(_GEN_21314); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21316 = 12'h824 == _T_643 ? $signed(7'sh26) : $signed(_GEN_21315); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21317 = 12'h825 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21316); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21318 = 12'h826 == _T_643 ? $signed(7'sh25) : $signed(_GEN_21317); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21319 = 12'h827 == _T_643 ? $signed(7'sh24) : $signed(_GEN_21318); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21320 = 12'h828 == _T_643 ? $signed(7'sh23) : $signed(_GEN_21319); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21321 = 12'h829 == _T_643 ? $signed(7'sh22) : $signed(_GEN_21320); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21322 = 12'h82a == _T_643 ? $signed(7'sh22) : $signed(_GEN_21321); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21323 = 12'h82b == _T_643 ? $signed(7'sh21) : $signed(_GEN_21322); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21324 = 12'h82c == _T_643 ? $signed(7'sh20) : $signed(_GEN_21323); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21325 = 12'h82d == _T_643 ? $signed(7'sh20) : $signed(_GEN_21324); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21326 = 12'h82e == _T_643 ? $signed(7'sh1f) : $signed(_GEN_21325); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21327 = 12'h82f == _T_643 ? $signed(7'sh1e) : $signed(_GEN_21326); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21328 = 12'h830 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21327); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21329 = 12'h831 == _T_643 ? $signed(7'sh1d) : $signed(_GEN_21328); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21330 = 12'h832 == _T_643 ? $signed(7'sh1c) : $signed(_GEN_21329); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21331 = 12'h833 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21330); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21332 = 12'h834 == _T_643 ? $signed(7'sh1b) : $signed(_GEN_21331); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21333 = 12'h835 == _T_643 ? $signed(7'sh1a) : $signed(_GEN_21332); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21334 = 12'h836 == _T_643 ? $signed(7'sh19) : $signed(_GEN_21333); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21335 = 12'h837 == _T_643 ? $signed(7'sh18) : $signed(_GEN_21334); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21336 = 12'h838 == _T_643 ? $signed(7'sh18) : $signed(_GEN_21335); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21337 = 12'h839 == _T_643 ? $signed(7'sh17) : $signed(_GEN_21336); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21338 = 12'h83a == _T_643 ? $signed(7'sh16) : $signed(_GEN_21337); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21339 = 12'h83b == _T_643 ? $signed(7'sh16) : $signed(_GEN_21338); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21340 = 12'h83c == _T_643 ? $signed(7'sh15) : $signed(_GEN_21339); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21341 = 12'h83d == _T_643 ? $signed(7'sh14) : $signed(_GEN_21340); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21342 = 12'h83e == _T_643 ? $signed(7'sh14) : $signed(_GEN_21341); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21343 = 12'h83f == _T_643 ? $signed(7'sh13) : $signed(_GEN_21342); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21344 = 12'h840 == _T_643 ? $signed(7'sh12) : $signed(_GEN_21343); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21345 = 12'h841 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21344); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21346 = 12'h842 == _T_643 ? $signed(7'sh11) : $signed(_GEN_21345); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_21347 = 12'h843 == _T_643 ? $signed(7'sh10) : $signed(_GEN_21346); // @[GraphicEngineVGA.scala 322:24]
  wire [11:0] _T_645 = spriteRotationReg_4 ? $signed({{5{_GEN_21347[6]}},_GEN_21347}) : $signed(_T_638); // @[GraphicEngineVGA.scala 322:24]
  wire  _T_646 = 2'h2 == spriteScaleHorizontalReg_4; // @[Mux.scala 80:60]
  wire [7:0] _T_647 = _T_646 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_648 = 2'h1 == spriteScaleHorizontalReg_4; // @[Mux.scala 80:60]
  wire [7:0] _T_649 = _T_648 ? $signed(8'sh10) : $signed(_T_647); // @[Mux.scala 80:57]
  wire  _T_650 = 2'h0 == spriteScaleHorizontalReg_4; // @[Mux.scala 80:60]
  wire [7:0] _T_651 = _T_650 ? $signed(8'sh20) : $signed(_T_649); // @[Mux.scala 80:57]
  wire  _T_652 = 2'h2 == spriteScaleVerticalReg_4; // @[Mux.scala 80:60]
  wire [7:0] _T_653 = _T_652 ? $signed(8'sh40) : $signed(8'sh20); // @[Mux.scala 80:57]
  wire  _T_654 = 2'h1 == spriteScaleVerticalReg_4; // @[Mux.scala 80:60]
  wire [7:0] _T_655 = _T_654 ? $signed(8'sh10) : $signed(_T_653); // @[Mux.scala 80:57]
  wire  _T_656 = 2'h0 == spriteScaleVerticalReg_4; // @[Mux.scala 80:60]
  wire [7:0] _T_657 = _T_656 ? $signed(8'sh20) : $signed(_T_655); // @[Mux.scala 80:57]
  wire [7:0] _T_660 = $signed(_T_651) - 8'sh1; // @[GraphicEngineVGA.scala 338:58]
  wire [11:0] _GEN_68002 = {{4{_T_660[7]}},_T_660}; // @[GraphicEngineVGA.scala 338:65]
  wire [11:0] _T_663 = $signed(_GEN_68002) - $signed(inSpriteX_4); // @[GraphicEngineVGA.scala 338:65]
  wire [11:0] _T_664 = spriteFlipHorizontalReg_4 ? $signed(_T_663) : $signed(inSpriteX_4); // @[GraphicEngineVGA.scala 338:23]
  wire [10:0] inSpriteY_4 = _T_645[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire  _T_672 = $signed(_T_628) >= 12'sh0; // @[GraphicEngineVGA.scala 343:27]
  wire  _T_673 = $signed(_T_628) < 12'sh2e; // @[GraphicEngineVGA.scala 343:47]
  wire  _T_674 = _T_672 & _T_673; // @[GraphicEngineVGA.scala 343:35]
  wire  _T_675 = $signed(_T_638) >= 12'sh0; // @[GraphicEngineVGA.scala 344:27]
  wire  _T_676 = $signed(_T_638) < 12'sh2e; // @[GraphicEngineVGA.scala 344:47]
  wire  _T_677 = _T_675 & _T_676; // @[GraphicEngineVGA.scala 344:35]
  wire  _T_678 = _T_674 & _T_677; // @[GraphicEngineVGA.scala 345:32]
  wire  _T_679 = $signed(_T_664) >= 12'sh0; // @[GraphicEngineVGA.scala 347:31]
  wire [11:0] _GEN_68005 = {{4{_T_651[7]}},_T_651}; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_680 = $signed(_T_664) < $signed(_GEN_68005); // @[GraphicEngineVGA.scala 347:52]
  wire  _T_681 = _T_679 & _T_680; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_682 = $signed(inSpriteY_4) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire [10:0] _GEN_68006 = {{3{_T_657[7]}},_T_657}; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_683 = $signed(inSpriteY_4) < $signed(_GEN_68006); // @[GraphicEngineVGA.scala 348:52]
  wire  _T_684 = _T_682 & _T_683; // @[GraphicEngineVGA.scala 348:39]
  wire  _T_685 = _T_678 & _T_681; // @[GraphicEngineVGA.scala 350:59]
  wire  _T_686 = _T_685 & _T_684; // @[GraphicEngineVGA.scala 350:72]
  wire  _T_687 = _T_681 & _T_684; // @[GraphicEngineVGA.scala 350:97]
  wire [10:0] _T_690 = _T_664[11:1]; // @[GraphicEngineVGA.scala 354:24]
  wire [6:0] _T_693 = _T_664[4:0] * 5'h2; // @[GraphicEngineVGA.scala 355:36]
  wire [4:0] _T_696 = _T_646 ? _T_690[4:0] : _T_664[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_698 = _T_648 ? _T_693 : {{2'd0}, _T_696}; // @[Mux.scala 80:57]
  wire [6:0] _T_700 = _T_650 ? {{2'd0}, _T_664[4:0]} : _T_698; // @[Mux.scala 80:57]
  wire [9:0] _T_702 = inSpriteY_4[10:1]; // @[GraphicEngineVGA.scala 359:24]
  wire [6:0] _T_705 = inSpriteY_4[4:0] * 5'h2; // @[GraphicEngineVGA.scala 360:36]
  wire [4:0] _T_708 = _T_652 ? _T_702[4:0] : inSpriteY_4[4:0]; // @[Mux.scala 80:57]
  wire [6:0] _T_710 = _T_654 ? _T_705 : {{2'd0}, _T_708}; // @[Mux.scala 80:57]
  wire [6:0] _T_712 = _T_656 ? {{2'd0}, inSpriteY_4[4:0]} : _T_710; // @[Mux.scala 80:57]
  wire [12:0] _T_713 = 7'h20 * _T_712; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_68007 = {{6'd0}, _T_700}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_715 = _GEN_68007 + _T_713; // @[GraphicEngineVGA.scala 367:46]
  wire [11:0] _T_718 = $signed(_T_232) - $signed(spriteXPositionReg_5); // @[GraphicEngineVGA.scala 301:73]
  wire [10:0] _GEN_68008 = {{1{spriteYPositionReg_5[9]}},spriteYPositionReg_5}; // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_728 = $signed(_T_242) - $signed(_GEN_68008); // @[GraphicEngineVGA.scala 302:73]
  wire [10:0] inSpriteY_5 = _T_728[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire [10:0] _T_767 = $signed(_GEN_67997) - $signed(inSpriteY_5); // @[GraphicEngineVGA.scala 339:65]
  wire [10:0] _T_768 = spriteFlipVerticalReg_5 ? $signed(_T_767) : $signed(inSpriteY_5); // @[GraphicEngineVGA.scala 339:23]
  wire  _T_769 = $signed(_T_718) >= 12'sh0; // @[GraphicEngineVGA.scala 343:27]
  wire  _T_777 = $signed(_T_718) < 12'sh20; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_778 = _T_769 & _T_777; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_779 = $signed(_T_768) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire  _T_780 = $signed(_T_768) < 11'sh20; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_781 = _T_779 & _T_780; // @[GraphicEngineVGA.scala 348:39]
  wire [6:0] _T_795 = {{2'd0}, _T_718[4:0]}; // @[Mux.scala 80:57]
  wire [6:0] _T_807 = {{2'd0}, _T_768[4:0]}; // @[Mux.scala 80:57]
  wire [12:0] _T_810 = 7'h20 * _T_807; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_68014 = {{6'd0}, _T_795}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_812 = _GEN_68014 + _T_810; // @[GraphicEngineVGA.scala 367:46]
  wire [11:0] _T_815 = $signed(_T_232) - $signed(spriteXPositionReg_6); // @[GraphicEngineVGA.scala 301:73]
  wire [11:0] _T_818 = $signed(_T_815) + 12'sh7; // @[GraphicEngineVGA.scala 301:98]
  wire [11:0] _T_822 = spriteRotationReg_6 ? $signed(_T_818) : $signed(_T_815); // @[GraphicEngineVGA.scala 301:22]
  wire [10:0] _GEN_68015 = {{1{spriteYPositionReg_6[9]}},spriteYPositionReg_6}; // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_825 = $signed(_T_242) - $signed(_GEN_68015); // @[GraphicEngineVGA.scala 302:73]
  wire [11:0] _T_828 = $signed(_T_825) + 12'sh7; // @[GraphicEngineVGA.scala 302:98]
  wire [11:0] _T_832 = spriteRotationReg_6 ? $signed(_T_828) : $signed(_T_825); // @[GraphicEngineVGA.scala 302:22]
  wire [11:0] _T_834 = _T_832[5:0] * 6'h2e; // @[GraphicEngineVGA.scala 307:34]
  wire [11:0] _GEN_68017 = {{6'd0}, _T_822[5:0]}; // @[GraphicEngineVGA.scala 307:53]
  wire [11:0] _T_837 = _T_834 + _GEN_68017; // @[GraphicEngineVGA.scala 307:53]
  wire [6:0] _GEN_25581 = 12'h1 == _T_837 ? $signed(-7'sh10) : $signed(-7'sh11); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25582 = 12'h2 == _T_837 ? $signed(-7'shf) : $signed(_GEN_25581); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25583 = 12'h3 == _T_837 ? $signed(-7'she) : $signed(_GEN_25582); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25584 = 12'h4 == _T_837 ? $signed(-7'she) : $signed(_GEN_25583); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25585 = 12'h5 == _T_837 ? $signed(-7'shd) : $signed(_GEN_25584); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25586 = 12'h6 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25585); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25587 = 12'h7 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25586); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25588 = 12'h8 == _T_837 ? $signed(-7'shb) : $signed(_GEN_25587); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25589 = 12'h9 == _T_837 ? $signed(-7'sha) : $signed(_GEN_25588); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25590 = 12'ha == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25589); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25591 = 12'hb == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25590); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25592 = 12'hc == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25591); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25593 = 12'hd == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25592); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25594 = 12'he == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25593); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25595 = 12'hf == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25594); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25596 = 12'h10 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25595); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25597 = 12'h11 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25596); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25598 = 12'h12 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25597); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25599 = 12'h13 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25598); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25600 = 12'h14 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25599); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25601 = 12'h15 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25600); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25602 = 12'h16 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25601); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25603 = 12'h17 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25602); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25604 = 12'h18 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25603); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25605 = 12'h19 == _T_837 ? $signed(7'sh1) : $signed(_GEN_25604); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25606 = 12'h1a == _T_837 ? $signed(7'sh2) : $signed(_GEN_25605); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25607 = 12'h1b == _T_837 ? $signed(7'sh3) : $signed(_GEN_25606); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25608 = 12'h1c == _T_837 ? $signed(7'sh3) : $signed(_GEN_25607); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25609 = 12'h1d == _T_837 ? $signed(7'sh4) : $signed(_GEN_25608); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25610 = 12'h1e == _T_837 ? $signed(7'sh5) : $signed(_GEN_25609); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25611 = 12'h1f == _T_837 ? $signed(7'sh5) : $signed(_GEN_25610); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25612 = 12'h20 == _T_837 ? $signed(7'sh6) : $signed(_GEN_25611); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25613 = 12'h21 == _T_837 ? $signed(7'sh7) : $signed(_GEN_25612); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25614 = 12'h22 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25613); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25615 = 12'h23 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25614); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25616 = 12'h24 == _T_837 ? $signed(7'sh9) : $signed(_GEN_25615); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25617 = 12'h25 == _T_837 ? $signed(7'sha) : $signed(_GEN_25616); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25618 = 12'h26 == _T_837 ? $signed(7'sha) : $signed(_GEN_25617); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25619 = 12'h27 == _T_837 ? $signed(7'shb) : $signed(_GEN_25618); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25620 = 12'h28 == _T_837 ? $signed(7'shc) : $signed(_GEN_25619); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25621 = 12'h29 == _T_837 ? $signed(7'shc) : $signed(_GEN_25620); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25622 = 12'h2a == _T_837 ? $signed(7'shd) : $signed(_GEN_25621); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25623 = 12'h2b == _T_837 ? $signed(7'she) : $signed(_GEN_25622); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25624 = 12'h2c == _T_837 ? $signed(7'shf) : $signed(_GEN_25623); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25625 = 12'h2d == _T_837 ? $signed(7'shf) : $signed(_GEN_25624); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25626 = 12'h2e == _T_837 ? $signed(-7'sh10) : $signed(_GEN_25625); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25627 = 12'h2f == _T_837 ? $signed(-7'shf) : $signed(_GEN_25626); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25628 = 12'h30 == _T_837 ? $signed(-7'she) : $signed(_GEN_25627); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25629 = 12'h31 == _T_837 ? $signed(-7'she) : $signed(_GEN_25628); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25630 = 12'h32 == _T_837 ? $signed(-7'shd) : $signed(_GEN_25629); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25631 = 12'h33 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25630); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25632 = 12'h34 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25631); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25633 = 12'h35 == _T_837 ? $signed(-7'shb) : $signed(_GEN_25632); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25634 = 12'h36 == _T_837 ? $signed(-7'sha) : $signed(_GEN_25633); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25635 = 12'h37 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25634); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25636 = 12'h38 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25635); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25637 = 12'h39 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25636); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25638 = 12'h3a == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25637); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25639 = 12'h3b == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25638); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25640 = 12'h3c == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25639); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25641 = 12'h3d == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25640); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25642 = 12'h3e == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25641); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25643 = 12'h3f == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25642); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25644 = 12'h40 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25643); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25645 = 12'h41 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25644); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25646 = 12'h42 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25645); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25647 = 12'h43 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25646); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25648 = 12'h44 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25647); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25649 = 12'h45 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25648); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25650 = 12'h46 == _T_837 ? $signed(7'sh1) : $signed(_GEN_25649); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25651 = 12'h47 == _T_837 ? $signed(7'sh2) : $signed(_GEN_25650); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25652 = 12'h48 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25651); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25653 = 12'h49 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25652); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25654 = 12'h4a == _T_837 ? $signed(7'sh4) : $signed(_GEN_25653); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25655 = 12'h4b == _T_837 ? $signed(7'sh5) : $signed(_GEN_25654); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25656 = 12'h4c == _T_837 ? $signed(7'sh5) : $signed(_GEN_25655); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25657 = 12'h4d == _T_837 ? $signed(7'sh6) : $signed(_GEN_25656); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25658 = 12'h4e == _T_837 ? $signed(7'sh7) : $signed(_GEN_25657); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25659 = 12'h4f == _T_837 ? $signed(7'sh8) : $signed(_GEN_25658); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25660 = 12'h50 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25659); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25661 = 12'h51 == _T_837 ? $signed(7'sh9) : $signed(_GEN_25660); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25662 = 12'h52 == _T_837 ? $signed(7'sha) : $signed(_GEN_25661); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25663 = 12'h53 == _T_837 ? $signed(7'sha) : $signed(_GEN_25662); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25664 = 12'h54 == _T_837 ? $signed(7'shb) : $signed(_GEN_25663); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25665 = 12'h55 == _T_837 ? $signed(7'shc) : $signed(_GEN_25664); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25666 = 12'h56 == _T_837 ? $signed(7'shc) : $signed(_GEN_25665); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25667 = 12'h57 == _T_837 ? $signed(7'shd) : $signed(_GEN_25666); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25668 = 12'h58 == _T_837 ? $signed(7'she) : $signed(_GEN_25667); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25669 = 12'h59 == _T_837 ? $signed(7'shf) : $signed(_GEN_25668); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25670 = 12'h5a == _T_837 ? $signed(7'shf) : $signed(_GEN_25669); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25671 = 12'h5b == _T_837 ? $signed(7'sh10) : $signed(_GEN_25670); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25672 = 12'h5c == _T_837 ? $signed(-7'shf) : $signed(_GEN_25671); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25673 = 12'h5d == _T_837 ? $signed(-7'she) : $signed(_GEN_25672); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25674 = 12'h5e == _T_837 ? $signed(-7'she) : $signed(_GEN_25673); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25675 = 12'h5f == _T_837 ? $signed(-7'shd) : $signed(_GEN_25674); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25676 = 12'h60 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25675); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25677 = 12'h61 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25676); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25678 = 12'h62 == _T_837 ? $signed(-7'shb) : $signed(_GEN_25677); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25679 = 12'h63 == _T_837 ? $signed(-7'sha) : $signed(_GEN_25678); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25680 = 12'h64 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25679); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25681 = 12'h65 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25680); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25682 = 12'h66 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25681); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25683 = 12'h67 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25682); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25684 = 12'h68 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25683); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25685 = 12'h69 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25684); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25686 = 12'h6a == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25685); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25687 = 12'h6b == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25686); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25688 = 12'h6c == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25687); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25689 = 12'h6d == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25688); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25690 = 12'h6e == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25689); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25691 = 12'h6f == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25690); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25692 = 12'h70 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25691); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25693 = 12'h71 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25692); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25694 = 12'h72 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25693); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25695 = 12'h73 == _T_837 ? $signed(7'sh1) : $signed(_GEN_25694); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25696 = 12'h74 == _T_837 ? $signed(7'sh2) : $signed(_GEN_25695); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25697 = 12'h75 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25696); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25698 = 12'h76 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25697); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25699 = 12'h77 == _T_837 ? $signed(7'sh4) : $signed(_GEN_25698); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25700 = 12'h78 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25699); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25701 = 12'h79 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25700); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25702 = 12'h7a == _T_837 ? $signed(7'sh6) : $signed(_GEN_25701); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25703 = 12'h7b == _T_837 ? $signed(7'sh7) : $signed(_GEN_25702); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25704 = 12'h7c == _T_837 ? $signed(7'sh8) : $signed(_GEN_25703); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25705 = 12'h7d == _T_837 ? $signed(7'sh8) : $signed(_GEN_25704); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25706 = 12'h7e == _T_837 ? $signed(7'sh9) : $signed(_GEN_25705); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25707 = 12'h7f == _T_837 ? $signed(7'sha) : $signed(_GEN_25706); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25708 = 12'h80 == _T_837 ? $signed(7'sha) : $signed(_GEN_25707); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25709 = 12'h81 == _T_837 ? $signed(7'shb) : $signed(_GEN_25708); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25710 = 12'h82 == _T_837 ? $signed(7'shc) : $signed(_GEN_25709); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25711 = 12'h83 == _T_837 ? $signed(7'shc) : $signed(_GEN_25710); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25712 = 12'h84 == _T_837 ? $signed(7'shd) : $signed(_GEN_25711); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25713 = 12'h85 == _T_837 ? $signed(7'she) : $signed(_GEN_25712); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25714 = 12'h86 == _T_837 ? $signed(7'shf) : $signed(_GEN_25713); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25715 = 12'h87 == _T_837 ? $signed(7'shf) : $signed(_GEN_25714); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25716 = 12'h88 == _T_837 ? $signed(7'sh10) : $signed(_GEN_25715); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25717 = 12'h89 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25716); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25718 = 12'h8a == _T_837 ? $signed(-7'she) : $signed(_GEN_25717); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25719 = 12'h8b == _T_837 ? $signed(-7'she) : $signed(_GEN_25718); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25720 = 12'h8c == _T_837 ? $signed(-7'shd) : $signed(_GEN_25719); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25721 = 12'h8d == _T_837 ? $signed(-7'shc) : $signed(_GEN_25720); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25722 = 12'h8e == _T_837 ? $signed(-7'shc) : $signed(_GEN_25721); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25723 = 12'h8f == _T_837 ? $signed(-7'shb) : $signed(_GEN_25722); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25724 = 12'h90 == _T_837 ? $signed(-7'sha) : $signed(_GEN_25723); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25725 = 12'h91 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25724); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25726 = 12'h92 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25725); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25727 = 12'h93 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25726); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25728 = 12'h94 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25727); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25729 = 12'h95 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25728); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25730 = 12'h96 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25729); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25731 = 12'h97 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25730); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25732 = 12'h98 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25731); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25733 = 12'h99 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25732); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25734 = 12'h9a == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25733); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25735 = 12'h9b == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25734); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25736 = 12'h9c == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25735); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25737 = 12'h9d == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25736); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25738 = 12'h9e == _T_837 ? $signed(7'sh0) : $signed(_GEN_25737); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25739 = 12'h9f == _T_837 ? $signed(7'sh0) : $signed(_GEN_25738); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25740 = 12'ha0 == _T_837 ? $signed(7'sh1) : $signed(_GEN_25739); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25741 = 12'ha1 == _T_837 ? $signed(7'sh2) : $signed(_GEN_25740); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25742 = 12'ha2 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25741); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25743 = 12'ha3 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25742); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25744 = 12'ha4 == _T_837 ? $signed(7'sh4) : $signed(_GEN_25743); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25745 = 12'ha5 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25744); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25746 = 12'ha6 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25745); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25747 = 12'ha7 == _T_837 ? $signed(7'sh6) : $signed(_GEN_25746); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25748 = 12'ha8 == _T_837 ? $signed(7'sh7) : $signed(_GEN_25747); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25749 = 12'ha9 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25748); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25750 = 12'haa == _T_837 ? $signed(7'sh8) : $signed(_GEN_25749); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25751 = 12'hab == _T_837 ? $signed(7'sh9) : $signed(_GEN_25750); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25752 = 12'hac == _T_837 ? $signed(7'sha) : $signed(_GEN_25751); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25753 = 12'had == _T_837 ? $signed(7'sha) : $signed(_GEN_25752); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25754 = 12'hae == _T_837 ? $signed(7'shb) : $signed(_GEN_25753); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25755 = 12'haf == _T_837 ? $signed(7'shc) : $signed(_GEN_25754); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25756 = 12'hb0 == _T_837 ? $signed(7'shc) : $signed(_GEN_25755); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25757 = 12'hb1 == _T_837 ? $signed(7'shd) : $signed(_GEN_25756); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25758 = 12'hb2 == _T_837 ? $signed(7'she) : $signed(_GEN_25757); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25759 = 12'hb3 == _T_837 ? $signed(7'shf) : $signed(_GEN_25758); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25760 = 12'hb4 == _T_837 ? $signed(7'shf) : $signed(_GEN_25759); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25761 = 12'hb5 == _T_837 ? $signed(7'sh10) : $signed(_GEN_25760); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25762 = 12'hb6 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25761); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25763 = 12'hb7 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25762); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25764 = 12'hb8 == _T_837 ? $signed(-7'she) : $signed(_GEN_25763); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25765 = 12'hb9 == _T_837 ? $signed(-7'shd) : $signed(_GEN_25764); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25766 = 12'hba == _T_837 ? $signed(-7'shc) : $signed(_GEN_25765); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25767 = 12'hbb == _T_837 ? $signed(-7'shc) : $signed(_GEN_25766); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25768 = 12'hbc == _T_837 ? $signed(-7'shb) : $signed(_GEN_25767); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25769 = 12'hbd == _T_837 ? $signed(-7'sha) : $signed(_GEN_25768); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25770 = 12'hbe == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25769); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25771 = 12'hbf == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25770); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25772 = 12'hc0 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25771); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25773 = 12'hc1 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25772); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25774 = 12'hc2 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25773); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25775 = 12'hc3 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25774); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25776 = 12'hc4 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25775); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25777 = 12'hc5 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25776); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25778 = 12'hc6 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25777); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25779 = 12'hc7 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25778); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25780 = 12'hc8 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25779); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25781 = 12'hc9 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25780); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25782 = 12'hca == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25781); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25783 = 12'hcb == _T_837 ? $signed(7'sh0) : $signed(_GEN_25782); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25784 = 12'hcc == _T_837 ? $signed(7'sh0) : $signed(_GEN_25783); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25785 = 12'hcd == _T_837 ? $signed(7'sh1) : $signed(_GEN_25784); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25786 = 12'hce == _T_837 ? $signed(7'sh2) : $signed(_GEN_25785); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25787 = 12'hcf == _T_837 ? $signed(7'sh3) : $signed(_GEN_25786); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25788 = 12'hd0 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25787); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25789 = 12'hd1 == _T_837 ? $signed(7'sh4) : $signed(_GEN_25788); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25790 = 12'hd2 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25789); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25791 = 12'hd3 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25790); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25792 = 12'hd4 == _T_837 ? $signed(7'sh6) : $signed(_GEN_25791); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25793 = 12'hd5 == _T_837 ? $signed(7'sh7) : $signed(_GEN_25792); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25794 = 12'hd6 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25793); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25795 = 12'hd7 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25794); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25796 = 12'hd8 == _T_837 ? $signed(7'sh9) : $signed(_GEN_25795); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25797 = 12'hd9 == _T_837 ? $signed(7'sha) : $signed(_GEN_25796); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25798 = 12'hda == _T_837 ? $signed(7'sha) : $signed(_GEN_25797); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25799 = 12'hdb == _T_837 ? $signed(7'shb) : $signed(_GEN_25798); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25800 = 12'hdc == _T_837 ? $signed(7'shc) : $signed(_GEN_25799); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25801 = 12'hdd == _T_837 ? $signed(7'shc) : $signed(_GEN_25800); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25802 = 12'hde == _T_837 ? $signed(7'shd) : $signed(_GEN_25801); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25803 = 12'hdf == _T_837 ? $signed(7'she) : $signed(_GEN_25802); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25804 = 12'he0 == _T_837 ? $signed(7'shf) : $signed(_GEN_25803); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25805 = 12'he1 == _T_837 ? $signed(7'shf) : $signed(_GEN_25804); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25806 = 12'he2 == _T_837 ? $signed(7'sh10) : $signed(_GEN_25805); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25807 = 12'he3 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25806); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25808 = 12'he4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25807); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25809 = 12'he5 == _T_837 ? $signed(7'sh12) : $signed(_GEN_25808); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25810 = 12'he6 == _T_837 ? $signed(-7'shd) : $signed(_GEN_25809); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25811 = 12'he7 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25810); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25812 = 12'he8 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25811); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25813 = 12'he9 == _T_837 ? $signed(-7'shb) : $signed(_GEN_25812); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25814 = 12'hea == _T_837 ? $signed(-7'sha) : $signed(_GEN_25813); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25815 = 12'heb == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25814); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25816 = 12'hec == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25815); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25817 = 12'hed == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25816); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25818 = 12'hee == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25817); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25819 = 12'hef == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25818); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25820 = 12'hf0 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25819); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25821 = 12'hf1 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25820); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25822 = 12'hf2 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25821); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25823 = 12'hf3 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25822); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25824 = 12'hf4 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25823); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25825 = 12'hf5 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25824); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25826 = 12'hf6 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25825); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25827 = 12'hf7 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25826); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25828 = 12'hf8 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25827); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25829 = 12'hf9 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25828); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25830 = 12'hfa == _T_837 ? $signed(7'sh1) : $signed(_GEN_25829); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25831 = 12'hfb == _T_837 ? $signed(7'sh2) : $signed(_GEN_25830); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25832 = 12'hfc == _T_837 ? $signed(7'sh3) : $signed(_GEN_25831); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25833 = 12'hfd == _T_837 ? $signed(7'sh3) : $signed(_GEN_25832); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25834 = 12'hfe == _T_837 ? $signed(7'sh4) : $signed(_GEN_25833); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25835 = 12'hff == _T_837 ? $signed(7'sh5) : $signed(_GEN_25834); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25836 = 12'h100 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25835); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25837 = 12'h101 == _T_837 ? $signed(7'sh6) : $signed(_GEN_25836); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25838 = 12'h102 == _T_837 ? $signed(7'sh7) : $signed(_GEN_25837); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25839 = 12'h103 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25838); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25840 = 12'h104 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25839); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25841 = 12'h105 == _T_837 ? $signed(7'sh9) : $signed(_GEN_25840); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25842 = 12'h106 == _T_837 ? $signed(7'sha) : $signed(_GEN_25841); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25843 = 12'h107 == _T_837 ? $signed(7'sha) : $signed(_GEN_25842); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25844 = 12'h108 == _T_837 ? $signed(7'shb) : $signed(_GEN_25843); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25845 = 12'h109 == _T_837 ? $signed(7'shc) : $signed(_GEN_25844); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25846 = 12'h10a == _T_837 ? $signed(7'shc) : $signed(_GEN_25845); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25847 = 12'h10b == _T_837 ? $signed(7'shd) : $signed(_GEN_25846); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25848 = 12'h10c == _T_837 ? $signed(7'she) : $signed(_GEN_25847); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25849 = 12'h10d == _T_837 ? $signed(7'shf) : $signed(_GEN_25848); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25850 = 12'h10e == _T_837 ? $signed(7'shf) : $signed(_GEN_25849); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25851 = 12'h10f == _T_837 ? $signed(7'sh10) : $signed(_GEN_25850); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25852 = 12'h110 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25851); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25853 = 12'h111 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25852); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25854 = 12'h112 == _T_837 ? $signed(7'sh12) : $signed(_GEN_25853); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25855 = 12'h113 == _T_837 ? $signed(7'sh13) : $signed(_GEN_25854); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25856 = 12'h114 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25855); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25857 = 12'h115 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25856); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25858 = 12'h116 == _T_837 ? $signed(-7'shb) : $signed(_GEN_25857); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25859 = 12'h117 == _T_837 ? $signed(-7'sha) : $signed(_GEN_25858); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25860 = 12'h118 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25859); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25861 = 12'h119 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25860); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25862 = 12'h11a == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25861); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25863 = 12'h11b == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25862); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25864 = 12'h11c == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25863); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25865 = 12'h11d == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25864); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25866 = 12'h11e == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25865); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25867 = 12'h11f == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25866); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25868 = 12'h120 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25867); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25869 = 12'h121 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25868); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25870 = 12'h122 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25869); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25871 = 12'h123 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25870); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25872 = 12'h124 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25871); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25873 = 12'h125 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25872); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25874 = 12'h126 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25873); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25875 = 12'h127 == _T_837 ? $signed(7'sh1) : $signed(_GEN_25874); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25876 = 12'h128 == _T_837 ? $signed(7'sh2) : $signed(_GEN_25875); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25877 = 12'h129 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25876); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25878 = 12'h12a == _T_837 ? $signed(7'sh3) : $signed(_GEN_25877); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25879 = 12'h12b == _T_837 ? $signed(7'sh4) : $signed(_GEN_25878); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25880 = 12'h12c == _T_837 ? $signed(7'sh5) : $signed(_GEN_25879); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25881 = 12'h12d == _T_837 ? $signed(7'sh5) : $signed(_GEN_25880); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25882 = 12'h12e == _T_837 ? $signed(7'sh6) : $signed(_GEN_25881); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25883 = 12'h12f == _T_837 ? $signed(7'sh7) : $signed(_GEN_25882); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25884 = 12'h130 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25883); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25885 = 12'h131 == _T_837 ? $signed(7'sh8) : $signed(_GEN_25884); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25886 = 12'h132 == _T_837 ? $signed(7'sh9) : $signed(_GEN_25885); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25887 = 12'h133 == _T_837 ? $signed(7'sha) : $signed(_GEN_25886); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25888 = 12'h134 == _T_837 ? $signed(7'sha) : $signed(_GEN_25887); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25889 = 12'h135 == _T_837 ? $signed(7'shb) : $signed(_GEN_25888); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25890 = 12'h136 == _T_837 ? $signed(7'shc) : $signed(_GEN_25889); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25891 = 12'h137 == _T_837 ? $signed(7'shc) : $signed(_GEN_25890); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25892 = 12'h138 == _T_837 ? $signed(7'shd) : $signed(_GEN_25891); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25893 = 12'h139 == _T_837 ? $signed(7'she) : $signed(_GEN_25892); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25894 = 12'h13a == _T_837 ? $signed(7'shf) : $signed(_GEN_25893); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25895 = 12'h13b == _T_837 ? $signed(7'shf) : $signed(_GEN_25894); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25896 = 12'h13c == _T_837 ? $signed(7'sh10) : $signed(_GEN_25895); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25897 = 12'h13d == _T_837 ? $signed(7'sh11) : $signed(_GEN_25896); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25898 = 12'h13e == _T_837 ? $signed(7'sh11) : $signed(_GEN_25897); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25899 = 12'h13f == _T_837 ? $signed(7'sh12) : $signed(_GEN_25898); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25900 = 12'h140 == _T_837 ? $signed(7'sh13) : $signed(_GEN_25899); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25901 = 12'h141 == _T_837 ? $signed(7'sh14) : $signed(_GEN_25900); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25902 = 12'h142 == _T_837 ? $signed(-7'shc) : $signed(_GEN_25901); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25903 = 12'h143 == _T_837 ? $signed(-7'shb) : $signed(_GEN_25902); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25904 = 12'h144 == _T_837 ? $signed(-7'sha) : $signed(_GEN_25903); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25905 = 12'h145 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25904); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25906 = 12'h146 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25905); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25907 = 12'h147 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25906); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25908 = 12'h148 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25907); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25909 = 12'h149 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25908); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25910 = 12'h14a == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25909); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25911 = 12'h14b == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25910); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25912 = 12'h14c == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25911); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25913 = 12'h14d == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25912); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25914 = 12'h14e == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25913); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25915 = 12'h14f == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25914); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25916 = 12'h150 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25915); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25917 = 12'h151 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25916); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25918 = 12'h152 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25917); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25919 = 12'h153 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25918); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25920 = 12'h154 == _T_837 ? $signed(7'sh1) : $signed(_GEN_25919); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25921 = 12'h155 == _T_837 ? $signed(7'sh2) : $signed(_GEN_25920); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25922 = 12'h156 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25921); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25923 = 12'h157 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25922); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25924 = 12'h158 == _T_837 ? $signed(7'sh4) : $signed(_GEN_25923); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25925 = 12'h159 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25924); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25926 = 12'h15a == _T_837 ? $signed(7'sh5) : $signed(_GEN_25925); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25927 = 12'h15b == _T_837 ? $signed(7'sh6) : $signed(_GEN_25926); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25928 = 12'h15c == _T_837 ? $signed(7'sh7) : $signed(_GEN_25927); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25929 = 12'h15d == _T_837 ? $signed(7'sh8) : $signed(_GEN_25928); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25930 = 12'h15e == _T_837 ? $signed(7'sh8) : $signed(_GEN_25929); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25931 = 12'h15f == _T_837 ? $signed(7'sh9) : $signed(_GEN_25930); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25932 = 12'h160 == _T_837 ? $signed(7'sha) : $signed(_GEN_25931); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25933 = 12'h161 == _T_837 ? $signed(7'sha) : $signed(_GEN_25932); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25934 = 12'h162 == _T_837 ? $signed(7'shb) : $signed(_GEN_25933); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25935 = 12'h163 == _T_837 ? $signed(7'shc) : $signed(_GEN_25934); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25936 = 12'h164 == _T_837 ? $signed(7'shc) : $signed(_GEN_25935); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25937 = 12'h165 == _T_837 ? $signed(7'shd) : $signed(_GEN_25936); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25938 = 12'h166 == _T_837 ? $signed(7'she) : $signed(_GEN_25937); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25939 = 12'h167 == _T_837 ? $signed(7'shf) : $signed(_GEN_25938); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25940 = 12'h168 == _T_837 ? $signed(7'shf) : $signed(_GEN_25939); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25941 = 12'h169 == _T_837 ? $signed(7'sh10) : $signed(_GEN_25940); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25942 = 12'h16a == _T_837 ? $signed(7'sh11) : $signed(_GEN_25941); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25943 = 12'h16b == _T_837 ? $signed(7'sh11) : $signed(_GEN_25942); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25944 = 12'h16c == _T_837 ? $signed(7'sh12) : $signed(_GEN_25943); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25945 = 12'h16d == _T_837 ? $signed(7'sh13) : $signed(_GEN_25944); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25946 = 12'h16e == _T_837 ? $signed(7'sh14) : $signed(_GEN_25945); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25947 = 12'h16f == _T_837 ? $signed(7'sh14) : $signed(_GEN_25946); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25948 = 12'h170 == _T_837 ? $signed(-7'shb) : $signed(_GEN_25947); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25949 = 12'h171 == _T_837 ? $signed(-7'sha) : $signed(_GEN_25948); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25950 = 12'h172 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25949); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25951 = 12'h173 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25950); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25952 = 12'h174 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25951); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25953 = 12'h175 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25952); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25954 = 12'h176 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25953); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25955 = 12'h177 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25954); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25956 = 12'h178 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25955); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25957 = 12'h179 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_25956); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25958 = 12'h17a == _T_837 ? $signed(-7'sh4) : $signed(_GEN_25957); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25959 = 12'h17b == _T_837 ? $signed(-7'sh3) : $signed(_GEN_25958); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25960 = 12'h17c == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25959); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25961 = 12'h17d == _T_837 ? $signed(-7'sh2) : $signed(_GEN_25960); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25962 = 12'h17e == _T_837 ? $signed(-7'sh1) : $signed(_GEN_25961); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25963 = 12'h17f == _T_837 ? $signed(7'sh0) : $signed(_GEN_25962); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25964 = 12'h180 == _T_837 ? $signed(7'sh0) : $signed(_GEN_25963); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25965 = 12'h181 == _T_837 ? $signed(7'sh1) : $signed(_GEN_25964); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25966 = 12'h182 == _T_837 ? $signed(7'sh2) : $signed(_GEN_25965); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25967 = 12'h183 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25966); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25968 = 12'h184 == _T_837 ? $signed(7'sh3) : $signed(_GEN_25967); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25969 = 12'h185 == _T_837 ? $signed(7'sh4) : $signed(_GEN_25968); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25970 = 12'h186 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25969); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25971 = 12'h187 == _T_837 ? $signed(7'sh5) : $signed(_GEN_25970); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25972 = 12'h188 == _T_837 ? $signed(7'sh6) : $signed(_GEN_25971); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25973 = 12'h189 == _T_837 ? $signed(7'sh7) : $signed(_GEN_25972); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25974 = 12'h18a == _T_837 ? $signed(7'sh8) : $signed(_GEN_25973); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25975 = 12'h18b == _T_837 ? $signed(7'sh8) : $signed(_GEN_25974); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25976 = 12'h18c == _T_837 ? $signed(7'sh9) : $signed(_GEN_25975); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25977 = 12'h18d == _T_837 ? $signed(7'sha) : $signed(_GEN_25976); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25978 = 12'h18e == _T_837 ? $signed(7'sha) : $signed(_GEN_25977); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25979 = 12'h18f == _T_837 ? $signed(7'shb) : $signed(_GEN_25978); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25980 = 12'h190 == _T_837 ? $signed(7'shc) : $signed(_GEN_25979); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25981 = 12'h191 == _T_837 ? $signed(7'shc) : $signed(_GEN_25980); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25982 = 12'h192 == _T_837 ? $signed(7'shd) : $signed(_GEN_25981); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25983 = 12'h193 == _T_837 ? $signed(7'she) : $signed(_GEN_25982); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25984 = 12'h194 == _T_837 ? $signed(7'shf) : $signed(_GEN_25983); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25985 = 12'h195 == _T_837 ? $signed(7'shf) : $signed(_GEN_25984); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25986 = 12'h196 == _T_837 ? $signed(7'sh10) : $signed(_GEN_25985); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25987 = 12'h197 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25986); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25988 = 12'h198 == _T_837 ? $signed(7'sh11) : $signed(_GEN_25987); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25989 = 12'h199 == _T_837 ? $signed(7'sh12) : $signed(_GEN_25988); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25990 = 12'h19a == _T_837 ? $signed(7'sh13) : $signed(_GEN_25989); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25991 = 12'h19b == _T_837 ? $signed(7'sh14) : $signed(_GEN_25990); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25992 = 12'h19c == _T_837 ? $signed(7'sh14) : $signed(_GEN_25991); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25993 = 12'h19d == _T_837 ? $signed(7'sh15) : $signed(_GEN_25992); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25994 = 12'h19e == _T_837 ? $signed(-7'sha) : $signed(_GEN_25993); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25995 = 12'h19f == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25994); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25996 = 12'h1a0 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_25995); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25997 = 12'h1a1 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_25996); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25998 = 12'h1a2 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25997); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_25999 = 12'h1a3 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_25998); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26000 = 12'h1a4 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_25999); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26001 = 12'h1a5 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26000); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26002 = 12'h1a6 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26001); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26003 = 12'h1a7 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26002); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26004 = 12'h1a8 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26003); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26005 = 12'h1a9 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26004); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26006 = 12'h1aa == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26005); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26007 = 12'h1ab == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26006); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26008 = 12'h1ac == _T_837 ? $signed(7'sh0) : $signed(_GEN_26007); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26009 = 12'h1ad == _T_837 ? $signed(7'sh0) : $signed(_GEN_26008); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26010 = 12'h1ae == _T_837 ? $signed(7'sh1) : $signed(_GEN_26009); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26011 = 12'h1af == _T_837 ? $signed(7'sh2) : $signed(_GEN_26010); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26012 = 12'h1b0 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26011); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26013 = 12'h1b1 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26012); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26014 = 12'h1b2 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26013); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26015 = 12'h1b3 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26014); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26016 = 12'h1b4 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26015); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26017 = 12'h1b5 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26016); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26018 = 12'h1b6 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26017); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26019 = 12'h1b7 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26018); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26020 = 12'h1b8 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26019); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26021 = 12'h1b9 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26020); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26022 = 12'h1ba == _T_837 ? $signed(7'sha) : $signed(_GEN_26021); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26023 = 12'h1bb == _T_837 ? $signed(7'sha) : $signed(_GEN_26022); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26024 = 12'h1bc == _T_837 ? $signed(7'shb) : $signed(_GEN_26023); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26025 = 12'h1bd == _T_837 ? $signed(7'shc) : $signed(_GEN_26024); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26026 = 12'h1be == _T_837 ? $signed(7'shc) : $signed(_GEN_26025); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26027 = 12'h1bf == _T_837 ? $signed(7'shd) : $signed(_GEN_26026); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26028 = 12'h1c0 == _T_837 ? $signed(7'she) : $signed(_GEN_26027); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26029 = 12'h1c1 == _T_837 ? $signed(7'shf) : $signed(_GEN_26028); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26030 = 12'h1c2 == _T_837 ? $signed(7'shf) : $signed(_GEN_26029); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26031 = 12'h1c3 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26030); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26032 = 12'h1c4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26031); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26033 = 12'h1c5 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26032); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26034 = 12'h1c6 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26033); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26035 = 12'h1c7 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26034); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26036 = 12'h1c8 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26035); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26037 = 12'h1c9 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26036); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26038 = 12'h1ca == _T_837 ? $signed(7'sh15) : $signed(_GEN_26037); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26039 = 12'h1cb == _T_837 ? $signed(7'sh16) : $signed(_GEN_26038); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26040 = 12'h1cc == _T_837 ? $signed(-7'sh9) : $signed(_GEN_26039); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26041 = 12'h1cd == _T_837 ? $signed(-7'sh9) : $signed(_GEN_26040); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26042 = 12'h1ce == _T_837 ? $signed(-7'sh8) : $signed(_GEN_26041); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26043 = 12'h1cf == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26042); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26044 = 12'h1d0 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26043); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26045 = 12'h1d1 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_26044); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26046 = 12'h1d2 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26045); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26047 = 12'h1d3 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26046); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26048 = 12'h1d4 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26047); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26049 = 12'h1d5 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26048); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26050 = 12'h1d6 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26049); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26051 = 12'h1d7 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26050); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26052 = 12'h1d8 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26051); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26053 = 12'h1d9 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26052); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26054 = 12'h1da == _T_837 ? $signed(7'sh0) : $signed(_GEN_26053); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26055 = 12'h1db == _T_837 ? $signed(7'sh1) : $signed(_GEN_26054); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26056 = 12'h1dc == _T_837 ? $signed(7'sh2) : $signed(_GEN_26055); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26057 = 12'h1dd == _T_837 ? $signed(7'sh3) : $signed(_GEN_26056); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26058 = 12'h1de == _T_837 ? $signed(7'sh3) : $signed(_GEN_26057); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26059 = 12'h1df == _T_837 ? $signed(7'sh4) : $signed(_GEN_26058); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26060 = 12'h1e0 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26059); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26061 = 12'h1e1 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26060); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26062 = 12'h1e2 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26061); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26063 = 12'h1e3 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26062); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26064 = 12'h1e4 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26063); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26065 = 12'h1e5 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26064); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26066 = 12'h1e6 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26065); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26067 = 12'h1e7 == _T_837 ? $signed(7'sha) : $signed(_GEN_26066); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26068 = 12'h1e8 == _T_837 ? $signed(7'sha) : $signed(_GEN_26067); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26069 = 12'h1e9 == _T_837 ? $signed(7'shb) : $signed(_GEN_26068); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26070 = 12'h1ea == _T_837 ? $signed(7'shc) : $signed(_GEN_26069); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26071 = 12'h1eb == _T_837 ? $signed(7'shc) : $signed(_GEN_26070); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26072 = 12'h1ec == _T_837 ? $signed(7'shd) : $signed(_GEN_26071); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26073 = 12'h1ed == _T_837 ? $signed(7'she) : $signed(_GEN_26072); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26074 = 12'h1ee == _T_837 ? $signed(7'shf) : $signed(_GEN_26073); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26075 = 12'h1ef == _T_837 ? $signed(7'shf) : $signed(_GEN_26074); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26076 = 12'h1f0 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26075); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26077 = 12'h1f1 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26076); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26078 = 12'h1f2 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26077); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26079 = 12'h1f3 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26078); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26080 = 12'h1f4 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26079); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26081 = 12'h1f5 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26080); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26082 = 12'h1f6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26081); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26083 = 12'h1f7 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26082); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26084 = 12'h1f8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26083); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26085 = 12'h1f9 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26084); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26086 = 12'h1fa == _T_837 ? $signed(-7'sh9) : $signed(_GEN_26085); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26087 = 12'h1fb == _T_837 ? $signed(-7'sh8) : $signed(_GEN_26086); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26088 = 12'h1fc == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26087); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26089 = 12'h1fd == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26088); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26090 = 12'h1fe == _T_837 ? $signed(-7'sh6) : $signed(_GEN_26089); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26091 = 12'h1ff == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26090); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26092 = 12'h200 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26091); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26093 = 12'h201 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26092); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26094 = 12'h202 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26093); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26095 = 12'h203 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26094); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26096 = 12'h204 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26095); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26097 = 12'h205 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26096); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26098 = 12'h206 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26097); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26099 = 12'h207 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26098); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26100 = 12'h208 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26099); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26101 = 12'h209 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26100); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26102 = 12'h20a == _T_837 ? $signed(7'sh3) : $signed(_GEN_26101); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26103 = 12'h20b == _T_837 ? $signed(7'sh3) : $signed(_GEN_26102); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26104 = 12'h20c == _T_837 ? $signed(7'sh4) : $signed(_GEN_26103); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26105 = 12'h20d == _T_837 ? $signed(7'sh5) : $signed(_GEN_26104); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26106 = 12'h20e == _T_837 ? $signed(7'sh5) : $signed(_GEN_26105); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26107 = 12'h20f == _T_837 ? $signed(7'sh6) : $signed(_GEN_26106); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26108 = 12'h210 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26107); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26109 = 12'h211 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26108); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26110 = 12'h212 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26109); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26111 = 12'h213 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26110); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26112 = 12'h214 == _T_837 ? $signed(7'sha) : $signed(_GEN_26111); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26113 = 12'h215 == _T_837 ? $signed(7'sha) : $signed(_GEN_26112); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26114 = 12'h216 == _T_837 ? $signed(7'shb) : $signed(_GEN_26113); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26115 = 12'h217 == _T_837 ? $signed(7'shc) : $signed(_GEN_26114); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26116 = 12'h218 == _T_837 ? $signed(7'shc) : $signed(_GEN_26115); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26117 = 12'h219 == _T_837 ? $signed(7'shd) : $signed(_GEN_26116); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26118 = 12'h21a == _T_837 ? $signed(7'she) : $signed(_GEN_26117); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26119 = 12'h21b == _T_837 ? $signed(7'shf) : $signed(_GEN_26118); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26120 = 12'h21c == _T_837 ? $signed(7'shf) : $signed(_GEN_26119); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26121 = 12'h21d == _T_837 ? $signed(7'sh10) : $signed(_GEN_26120); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26122 = 12'h21e == _T_837 ? $signed(7'sh11) : $signed(_GEN_26121); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26123 = 12'h21f == _T_837 ? $signed(7'sh11) : $signed(_GEN_26122); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26124 = 12'h220 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26123); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26125 = 12'h221 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26124); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26126 = 12'h222 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26125); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26127 = 12'h223 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26126); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26128 = 12'h224 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26127); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26129 = 12'h225 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26128); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26130 = 12'h226 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26129); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26131 = 12'h227 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26130); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26132 = 12'h228 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_26131); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26133 = 12'h229 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26132); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26134 = 12'h22a == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26133); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26135 = 12'h22b == _T_837 ? $signed(-7'sh6) : $signed(_GEN_26134); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26136 = 12'h22c == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26135); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26137 = 12'h22d == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26136); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26138 = 12'h22e == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26137); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26139 = 12'h22f == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26138); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26140 = 12'h230 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26139); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26141 = 12'h231 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26140); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26142 = 12'h232 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26141); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26143 = 12'h233 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26142); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26144 = 12'h234 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26143); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26145 = 12'h235 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26144); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26146 = 12'h236 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26145); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26147 = 12'h237 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26146); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26148 = 12'h238 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26147); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26149 = 12'h239 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26148); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26150 = 12'h23a == _T_837 ? $signed(7'sh5) : $signed(_GEN_26149); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26151 = 12'h23b == _T_837 ? $signed(7'sh5) : $signed(_GEN_26150); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26152 = 12'h23c == _T_837 ? $signed(7'sh6) : $signed(_GEN_26151); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26153 = 12'h23d == _T_837 ? $signed(7'sh7) : $signed(_GEN_26152); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26154 = 12'h23e == _T_837 ? $signed(7'sh8) : $signed(_GEN_26153); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26155 = 12'h23f == _T_837 ? $signed(7'sh8) : $signed(_GEN_26154); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26156 = 12'h240 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26155); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26157 = 12'h241 == _T_837 ? $signed(7'sha) : $signed(_GEN_26156); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26158 = 12'h242 == _T_837 ? $signed(7'sha) : $signed(_GEN_26157); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26159 = 12'h243 == _T_837 ? $signed(7'shb) : $signed(_GEN_26158); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26160 = 12'h244 == _T_837 ? $signed(7'shc) : $signed(_GEN_26159); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26161 = 12'h245 == _T_837 ? $signed(7'shc) : $signed(_GEN_26160); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26162 = 12'h246 == _T_837 ? $signed(7'shd) : $signed(_GEN_26161); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26163 = 12'h247 == _T_837 ? $signed(7'she) : $signed(_GEN_26162); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26164 = 12'h248 == _T_837 ? $signed(7'shf) : $signed(_GEN_26163); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26165 = 12'h249 == _T_837 ? $signed(7'shf) : $signed(_GEN_26164); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26166 = 12'h24a == _T_837 ? $signed(7'sh10) : $signed(_GEN_26165); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26167 = 12'h24b == _T_837 ? $signed(7'sh11) : $signed(_GEN_26166); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26168 = 12'h24c == _T_837 ? $signed(7'sh11) : $signed(_GEN_26167); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26169 = 12'h24d == _T_837 ? $signed(7'sh12) : $signed(_GEN_26168); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26170 = 12'h24e == _T_837 ? $signed(7'sh13) : $signed(_GEN_26169); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26171 = 12'h24f == _T_837 ? $signed(7'sh14) : $signed(_GEN_26170); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26172 = 12'h250 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26171); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26173 = 12'h251 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26172); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26174 = 12'h252 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26173); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26175 = 12'h253 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26174); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26176 = 12'h254 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26175); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26177 = 12'h255 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26176); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26178 = 12'h256 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26177); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26179 = 12'h257 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26178); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26180 = 12'h258 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_26179); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26181 = 12'h259 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26180); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26182 = 12'h25a == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26181); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26183 = 12'h25b == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26182); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26184 = 12'h25c == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26183); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26185 = 12'h25d == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26184); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26186 = 12'h25e == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26185); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26187 = 12'h25f == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26186); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26188 = 12'h260 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26187); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26189 = 12'h261 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26188); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26190 = 12'h262 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26189); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26191 = 12'h263 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26190); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26192 = 12'h264 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26191); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26193 = 12'h265 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26192); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26194 = 12'h266 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26193); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26195 = 12'h267 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26194); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26196 = 12'h268 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26195); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26197 = 12'h269 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26196); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26198 = 12'h26a == _T_837 ? $signed(7'sh7) : $signed(_GEN_26197); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26199 = 12'h26b == _T_837 ? $signed(7'sh8) : $signed(_GEN_26198); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26200 = 12'h26c == _T_837 ? $signed(7'sh8) : $signed(_GEN_26199); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26201 = 12'h26d == _T_837 ? $signed(7'sh9) : $signed(_GEN_26200); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26202 = 12'h26e == _T_837 ? $signed(7'sha) : $signed(_GEN_26201); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26203 = 12'h26f == _T_837 ? $signed(7'sha) : $signed(_GEN_26202); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26204 = 12'h270 == _T_837 ? $signed(7'shb) : $signed(_GEN_26203); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26205 = 12'h271 == _T_837 ? $signed(7'shc) : $signed(_GEN_26204); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26206 = 12'h272 == _T_837 ? $signed(7'shc) : $signed(_GEN_26205); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26207 = 12'h273 == _T_837 ? $signed(7'shd) : $signed(_GEN_26206); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26208 = 12'h274 == _T_837 ? $signed(7'she) : $signed(_GEN_26207); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26209 = 12'h275 == _T_837 ? $signed(7'shf) : $signed(_GEN_26208); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26210 = 12'h276 == _T_837 ? $signed(7'shf) : $signed(_GEN_26209); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26211 = 12'h277 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26210); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26212 = 12'h278 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26211); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26213 = 12'h279 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26212); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26214 = 12'h27a == _T_837 ? $signed(7'sh12) : $signed(_GEN_26213); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26215 = 12'h27b == _T_837 ? $signed(7'sh13) : $signed(_GEN_26214); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26216 = 12'h27c == _T_837 ? $signed(7'sh14) : $signed(_GEN_26215); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26217 = 12'h27d == _T_837 ? $signed(7'sh14) : $signed(_GEN_26216); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26218 = 12'h27e == _T_837 ? $signed(7'sh15) : $signed(_GEN_26217); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26219 = 12'h27f == _T_837 ? $signed(7'sh16) : $signed(_GEN_26218); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26220 = 12'h280 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26219); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26221 = 12'h281 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26220); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26222 = 12'h282 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26221); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26223 = 12'h283 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26222); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26224 = 12'h284 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_26223); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26225 = 12'h285 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_26224); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26226 = 12'h286 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26225); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26227 = 12'h287 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26226); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26228 = 12'h288 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26227); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26229 = 12'h289 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26228); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26230 = 12'h28a == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26229); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26231 = 12'h28b == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26230); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26232 = 12'h28c == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26231); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26233 = 12'h28d == _T_837 ? $signed(7'sh0) : $signed(_GEN_26232); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26234 = 12'h28e == _T_837 ? $signed(7'sh0) : $signed(_GEN_26233); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26235 = 12'h28f == _T_837 ? $signed(7'sh1) : $signed(_GEN_26234); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26236 = 12'h290 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26235); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26237 = 12'h291 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26236); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26238 = 12'h292 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26237); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26239 = 12'h293 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26238); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26240 = 12'h294 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26239); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26241 = 12'h295 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26240); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26242 = 12'h296 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26241); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26243 = 12'h297 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26242); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26244 = 12'h298 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26243); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26245 = 12'h299 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26244); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26246 = 12'h29a == _T_837 ? $signed(7'sh9) : $signed(_GEN_26245); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26247 = 12'h29b == _T_837 ? $signed(7'sha) : $signed(_GEN_26246); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26248 = 12'h29c == _T_837 ? $signed(7'sha) : $signed(_GEN_26247); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26249 = 12'h29d == _T_837 ? $signed(7'shb) : $signed(_GEN_26248); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26250 = 12'h29e == _T_837 ? $signed(7'shc) : $signed(_GEN_26249); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26251 = 12'h29f == _T_837 ? $signed(7'shc) : $signed(_GEN_26250); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26252 = 12'h2a0 == _T_837 ? $signed(7'shd) : $signed(_GEN_26251); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26253 = 12'h2a1 == _T_837 ? $signed(7'she) : $signed(_GEN_26252); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26254 = 12'h2a2 == _T_837 ? $signed(7'shf) : $signed(_GEN_26253); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26255 = 12'h2a3 == _T_837 ? $signed(7'shf) : $signed(_GEN_26254); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26256 = 12'h2a4 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26255); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26257 = 12'h2a5 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26256); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26258 = 12'h2a6 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26257); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26259 = 12'h2a7 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26258); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26260 = 12'h2a8 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26259); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26261 = 12'h2a9 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26260); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26262 = 12'h2aa == _T_837 ? $signed(7'sh14) : $signed(_GEN_26261); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26263 = 12'h2ab == _T_837 ? $signed(7'sh15) : $signed(_GEN_26262); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26264 = 12'h2ac == _T_837 ? $signed(7'sh16) : $signed(_GEN_26263); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26265 = 12'h2ad == _T_837 ? $signed(7'sh16) : $signed(_GEN_26264); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26266 = 12'h2ae == _T_837 ? $signed(7'sh17) : $signed(_GEN_26265); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26267 = 12'h2af == _T_837 ? $signed(7'sh18) : $signed(_GEN_26266); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26268 = 12'h2b0 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26267); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26269 = 12'h2b1 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26268); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26270 = 12'h2b2 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_26269); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26271 = 12'h2b3 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26270); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26272 = 12'h2b4 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26271); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26273 = 12'h2b5 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26272); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26274 = 12'h2b6 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26273); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26275 = 12'h2b7 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26274); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26276 = 12'h2b8 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26275); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26277 = 12'h2b9 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26276); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26278 = 12'h2ba == _T_837 ? $signed(7'sh0) : $signed(_GEN_26277); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26279 = 12'h2bb == _T_837 ? $signed(7'sh0) : $signed(_GEN_26278); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26280 = 12'h2bc == _T_837 ? $signed(7'sh1) : $signed(_GEN_26279); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26281 = 12'h2bd == _T_837 ? $signed(7'sh2) : $signed(_GEN_26280); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26282 = 12'h2be == _T_837 ? $signed(7'sh3) : $signed(_GEN_26281); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26283 = 12'h2bf == _T_837 ? $signed(7'sh3) : $signed(_GEN_26282); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26284 = 12'h2c0 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26283); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26285 = 12'h2c1 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26284); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26286 = 12'h2c2 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26285); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26287 = 12'h2c3 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26286); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26288 = 12'h2c4 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26287); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26289 = 12'h2c5 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26288); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26290 = 12'h2c6 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26289); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26291 = 12'h2c7 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26290); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26292 = 12'h2c8 == _T_837 ? $signed(7'sha) : $signed(_GEN_26291); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26293 = 12'h2c9 == _T_837 ? $signed(7'sha) : $signed(_GEN_26292); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26294 = 12'h2ca == _T_837 ? $signed(7'shb) : $signed(_GEN_26293); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26295 = 12'h2cb == _T_837 ? $signed(7'shc) : $signed(_GEN_26294); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26296 = 12'h2cc == _T_837 ? $signed(7'shc) : $signed(_GEN_26295); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26297 = 12'h2cd == _T_837 ? $signed(7'shd) : $signed(_GEN_26296); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26298 = 12'h2ce == _T_837 ? $signed(7'she) : $signed(_GEN_26297); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26299 = 12'h2cf == _T_837 ? $signed(7'shf) : $signed(_GEN_26298); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26300 = 12'h2d0 == _T_837 ? $signed(7'shf) : $signed(_GEN_26299); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26301 = 12'h2d1 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26300); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26302 = 12'h2d2 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26301); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26303 = 12'h2d3 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26302); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26304 = 12'h2d4 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26303); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26305 = 12'h2d5 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26304); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26306 = 12'h2d6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26305); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26307 = 12'h2d7 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26306); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26308 = 12'h2d8 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26307); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26309 = 12'h2d9 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26308); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26310 = 12'h2da == _T_837 ? $signed(7'sh16) : $signed(_GEN_26309); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26311 = 12'h2db == _T_837 ? $signed(7'sh17) : $signed(_GEN_26310); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26312 = 12'h2dc == _T_837 ? $signed(7'sh18) : $signed(_GEN_26311); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26313 = 12'h2dd == _T_837 ? $signed(7'sh18) : $signed(_GEN_26312); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26314 = 12'h2de == _T_837 ? $signed(7'sh19) : $signed(_GEN_26313); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26315 = 12'h2df == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26314); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26316 = 12'h2e0 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26315); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26317 = 12'h2e1 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26316); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26318 = 12'h2e2 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26317); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26319 = 12'h2e3 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26318); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26320 = 12'h2e4 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26319); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26321 = 12'h2e5 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26320); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26322 = 12'h2e6 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26321); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26323 = 12'h2e7 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26322); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26324 = 12'h2e8 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26323); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26325 = 12'h2e9 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26324); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26326 = 12'h2ea == _T_837 ? $signed(7'sh2) : $signed(_GEN_26325); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26327 = 12'h2eb == _T_837 ? $signed(7'sh3) : $signed(_GEN_26326); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26328 = 12'h2ec == _T_837 ? $signed(7'sh3) : $signed(_GEN_26327); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26329 = 12'h2ed == _T_837 ? $signed(7'sh4) : $signed(_GEN_26328); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26330 = 12'h2ee == _T_837 ? $signed(7'sh5) : $signed(_GEN_26329); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26331 = 12'h2ef == _T_837 ? $signed(7'sh5) : $signed(_GEN_26330); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26332 = 12'h2f0 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26331); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26333 = 12'h2f1 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26332); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26334 = 12'h2f2 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26333); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26335 = 12'h2f3 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26334); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26336 = 12'h2f4 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26335); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26337 = 12'h2f5 == _T_837 ? $signed(7'sha) : $signed(_GEN_26336); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26338 = 12'h2f6 == _T_837 ? $signed(7'sha) : $signed(_GEN_26337); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26339 = 12'h2f7 == _T_837 ? $signed(7'shb) : $signed(_GEN_26338); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26340 = 12'h2f8 == _T_837 ? $signed(7'shc) : $signed(_GEN_26339); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26341 = 12'h2f9 == _T_837 ? $signed(7'shc) : $signed(_GEN_26340); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26342 = 12'h2fa == _T_837 ? $signed(7'shd) : $signed(_GEN_26341); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26343 = 12'h2fb == _T_837 ? $signed(7'she) : $signed(_GEN_26342); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26344 = 12'h2fc == _T_837 ? $signed(7'shf) : $signed(_GEN_26343); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26345 = 12'h2fd == _T_837 ? $signed(7'shf) : $signed(_GEN_26344); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26346 = 12'h2fe == _T_837 ? $signed(7'sh10) : $signed(_GEN_26345); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26347 = 12'h2ff == _T_837 ? $signed(7'sh11) : $signed(_GEN_26346); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26348 = 12'h300 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26347); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26349 = 12'h301 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26348); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26350 = 12'h302 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26349); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26351 = 12'h303 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26350); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26352 = 12'h304 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26351); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26353 = 12'h305 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26352); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26354 = 12'h306 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26353); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26355 = 12'h307 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26354); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26356 = 12'h308 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26355); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26357 = 12'h309 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26356); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26358 = 12'h30a == _T_837 ? $signed(7'sh18) : $signed(_GEN_26357); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26359 = 12'h30b == _T_837 ? $signed(7'sh19) : $signed(_GEN_26358); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26360 = 12'h30c == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26359); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26361 = 12'h30d == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26360); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26362 = 12'h30e == _T_837 ? $signed(-7'sh5) : $signed(_GEN_26361); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26363 = 12'h30f == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26362); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26364 = 12'h310 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26363); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26365 = 12'h311 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26364); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26366 = 12'h312 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26365); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26367 = 12'h313 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26366); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26368 = 12'h314 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26367); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26369 = 12'h315 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26368); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26370 = 12'h316 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26369); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26371 = 12'h317 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26370); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26372 = 12'h318 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26371); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26373 = 12'h319 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26372); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26374 = 12'h31a == _T_837 ? $signed(7'sh4) : $signed(_GEN_26373); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26375 = 12'h31b == _T_837 ? $signed(7'sh5) : $signed(_GEN_26374); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26376 = 12'h31c == _T_837 ? $signed(7'sh5) : $signed(_GEN_26375); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26377 = 12'h31d == _T_837 ? $signed(7'sh6) : $signed(_GEN_26376); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26378 = 12'h31e == _T_837 ? $signed(7'sh7) : $signed(_GEN_26377); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26379 = 12'h31f == _T_837 ? $signed(7'sh8) : $signed(_GEN_26378); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26380 = 12'h320 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26379); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26381 = 12'h321 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26380); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26382 = 12'h322 == _T_837 ? $signed(7'sha) : $signed(_GEN_26381); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26383 = 12'h323 == _T_837 ? $signed(7'sha) : $signed(_GEN_26382); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26384 = 12'h324 == _T_837 ? $signed(7'shb) : $signed(_GEN_26383); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26385 = 12'h325 == _T_837 ? $signed(7'shc) : $signed(_GEN_26384); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26386 = 12'h326 == _T_837 ? $signed(7'shc) : $signed(_GEN_26385); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26387 = 12'h327 == _T_837 ? $signed(7'shd) : $signed(_GEN_26386); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26388 = 12'h328 == _T_837 ? $signed(7'she) : $signed(_GEN_26387); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26389 = 12'h329 == _T_837 ? $signed(7'shf) : $signed(_GEN_26388); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26390 = 12'h32a == _T_837 ? $signed(7'shf) : $signed(_GEN_26389); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26391 = 12'h32b == _T_837 ? $signed(7'sh10) : $signed(_GEN_26390); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26392 = 12'h32c == _T_837 ? $signed(7'sh11) : $signed(_GEN_26391); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26393 = 12'h32d == _T_837 ? $signed(7'sh11) : $signed(_GEN_26392); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26394 = 12'h32e == _T_837 ? $signed(7'sh12) : $signed(_GEN_26393); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26395 = 12'h32f == _T_837 ? $signed(7'sh13) : $signed(_GEN_26394); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26396 = 12'h330 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26395); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26397 = 12'h331 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26396); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26398 = 12'h332 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26397); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26399 = 12'h333 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26398); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26400 = 12'h334 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26399); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26401 = 12'h335 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26400); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26402 = 12'h336 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26401); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26403 = 12'h337 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26402); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26404 = 12'h338 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26403); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26405 = 12'h339 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26404); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26406 = 12'h33a == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26405); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26407 = 12'h33b == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26406); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26408 = 12'h33c == _T_837 ? $signed(-7'sh4) : $signed(_GEN_26407); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26409 = 12'h33d == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26408); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26410 = 12'h33e == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26409); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26411 = 12'h33f == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26410); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26412 = 12'h340 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26411); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26413 = 12'h341 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26412); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26414 = 12'h342 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26413); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26415 = 12'h343 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26414); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26416 = 12'h344 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26415); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26417 = 12'h345 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26416); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26418 = 12'h346 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26417); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26419 = 12'h347 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26418); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26420 = 12'h348 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26419); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26421 = 12'h349 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26420); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26422 = 12'h34a == _T_837 ? $signed(7'sh6) : $signed(_GEN_26421); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26423 = 12'h34b == _T_837 ? $signed(7'sh7) : $signed(_GEN_26422); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26424 = 12'h34c == _T_837 ? $signed(7'sh8) : $signed(_GEN_26423); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26425 = 12'h34d == _T_837 ? $signed(7'sh8) : $signed(_GEN_26424); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26426 = 12'h34e == _T_837 ? $signed(7'sh9) : $signed(_GEN_26425); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26427 = 12'h34f == _T_837 ? $signed(7'sha) : $signed(_GEN_26426); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26428 = 12'h350 == _T_837 ? $signed(7'sha) : $signed(_GEN_26427); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26429 = 12'h351 == _T_837 ? $signed(7'shb) : $signed(_GEN_26428); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26430 = 12'h352 == _T_837 ? $signed(7'shc) : $signed(_GEN_26429); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26431 = 12'h353 == _T_837 ? $signed(7'shc) : $signed(_GEN_26430); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26432 = 12'h354 == _T_837 ? $signed(7'shd) : $signed(_GEN_26431); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26433 = 12'h355 == _T_837 ? $signed(7'she) : $signed(_GEN_26432); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26434 = 12'h356 == _T_837 ? $signed(7'shf) : $signed(_GEN_26433); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26435 = 12'h357 == _T_837 ? $signed(7'shf) : $signed(_GEN_26434); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26436 = 12'h358 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26435); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26437 = 12'h359 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26436); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26438 = 12'h35a == _T_837 ? $signed(7'sh11) : $signed(_GEN_26437); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26439 = 12'h35b == _T_837 ? $signed(7'sh12) : $signed(_GEN_26438); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26440 = 12'h35c == _T_837 ? $signed(7'sh13) : $signed(_GEN_26439); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26441 = 12'h35d == _T_837 ? $signed(7'sh14) : $signed(_GEN_26440); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26442 = 12'h35e == _T_837 ? $signed(7'sh14) : $signed(_GEN_26441); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26443 = 12'h35f == _T_837 ? $signed(7'sh15) : $signed(_GEN_26442); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26444 = 12'h360 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26443); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26445 = 12'h361 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26444); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26446 = 12'h362 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26445); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26447 = 12'h363 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26446); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26448 = 12'h364 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26447); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26449 = 12'h365 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26448); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26450 = 12'h366 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26449); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26451 = 12'h367 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26450); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26452 = 12'h368 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26451); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26453 = 12'h369 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26452); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26454 = 12'h36a == _T_837 ? $signed(-7'sh3) : $signed(_GEN_26453); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26455 = 12'h36b == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26454); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26456 = 12'h36c == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26455); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26457 = 12'h36d == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26456); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26458 = 12'h36e == _T_837 ? $signed(7'sh0) : $signed(_GEN_26457); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26459 = 12'h36f == _T_837 ? $signed(7'sh0) : $signed(_GEN_26458); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26460 = 12'h370 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26459); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26461 = 12'h371 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26460); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26462 = 12'h372 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26461); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26463 = 12'h373 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26462); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26464 = 12'h374 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26463); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26465 = 12'h375 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26464); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26466 = 12'h376 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26465); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26467 = 12'h377 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26466); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26468 = 12'h378 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26467); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26469 = 12'h379 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26468); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26470 = 12'h37a == _T_837 ? $signed(7'sh8) : $signed(_GEN_26469); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26471 = 12'h37b == _T_837 ? $signed(7'sh9) : $signed(_GEN_26470); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26472 = 12'h37c == _T_837 ? $signed(7'sha) : $signed(_GEN_26471); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26473 = 12'h37d == _T_837 ? $signed(7'sha) : $signed(_GEN_26472); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26474 = 12'h37e == _T_837 ? $signed(7'shb) : $signed(_GEN_26473); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26475 = 12'h37f == _T_837 ? $signed(7'shc) : $signed(_GEN_26474); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26476 = 12'h380 == _T_837 ? $signed(7'shc) : $signed(_GEN_26475); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26477 = 12'h381 == _T_837 ? $signed(7'shd) : $signed(_GEN_26476); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26478 = 12'h382 == _T_837 ? $signed(7'she) : $signed(_GEN_26477); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26479 = 12'h383 == _T_837 ? $signed(7'shf) : $signed(_GEN_26478); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26480 = 12'h384 == _T_837 ? $signed(7'shf) : $signed(_GEN_26479); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26481 = 12'h385 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26480); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26482 = 12'h386 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26481); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26483 = 12'h387 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26482); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26484 = 12'h388 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26483); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26485 = 12'h389 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26484); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26486 = 12'h38a == _T_837 ? $signed(7'sh14) : $signed(_GEN_26485); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26487 = 12'h38b == _T_837 ? $signed(7'sh14) : $signed(_GEN_26486); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26488 = 12'h38c == _T_837 ? $signed(7'sh15) : $signed(_GEN_26487); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26489 = 12'h38d == _T_837 ? $signed(7'sh16) : $signed(_GEN_26488); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26490 = 12'h38e == _T_837 ? $signed(7'sh16) : $signed(_GEN_26489); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26491 = 12'h38f == _T_837 ? $signed(7'sh17) : $signed(_GEN_26490); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26492 = 12'h390 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26491); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26493 = 12'h391 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26492); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26494 = 12'h392 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26493); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26495 = 12'h393 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26494); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26496 = 12'h394 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26495); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26497 = 12'h395 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26496); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26498 = 12'h396 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26497); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26499 = 12'h397 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26498); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26500 = 12'h398 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26499); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26501 = 12'h399 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26500); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26502 = 12'h39a == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26501); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26503 = 12'h39b == _T_837 ? $signed(7'sh0) : $signed(_GEN_26502); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26504 = 12'h39c == _T_837 ? $signed(7'sh0) : $signed(_GEN_26503); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26505 = 12'h39d == _T_837 ? $signed(7'sh1) : $signed(_GEN_26504); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26506 = 12'h39e == _T_837 ? $signed(7'sh2) : $signed(_GEN_26505); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26507 = 12'h39f == _T_837 ? $signed(7'sh3) : $signed(_GEN_26506); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26508 = 12'h3a0 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26507); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26509 = 12'h3a1 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26508); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26510 = 12'h3a2 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26509); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26511 = 12'h3a3 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26510); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26512 = 12'h3a4 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26511); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26513 = 12'h3a5 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26512); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26514 = 12'h3a6 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26513); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26515 = 12'h3a7 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26514); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26516 = 12'h3a8 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26515); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26517 = 12'h3a9 == _T_837 ? $signed(7'sha) : $signed(_GEN_26516); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26518 = 12'h3aa == _T_837 ? $signed(7'sha) : $signed(_GEN_26517); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26519 = 12'h3ab == _T_837 ? $signed(7'shb) : $signed(_GEN_26518); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26520 = 12'h3ac == _T_837 ? $signed(7'shc) : $signed(_GEN_26519); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26521 = 12'h3ad == _T_837 ? $signed(7'shc) : $signed(_GEN_26520); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26522 = 12'h3ae == _T_837 ? $signed(7'shd) : $signed(_GEN_26521); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26523 = 12'h3af == _T_837 ? $signed(7'she) : $signed(_GEN_26522); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26524 = 12'h3b0 == _T_837 ? $signed(7'shf) : $signed(_GEN_26523); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26525 = 12'h3b1 == _T_837 ? $signed(7'shf) : $signed(_GEN_26524); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26526 = 12'h3b2 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26525); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26527 = 12'h3b3 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26526); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26528 = 12'h3b4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26527); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26529 = 12'h3b5 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26528); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26530 = 12'h3b6 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26529); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26531 = 12'h3b7 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26530); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26532 = 12'h3b8 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26531); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26533 = 12'h3b9 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26532); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26534 = 12'h3ba == _T_837 ? $signed(7'sh16) : $signed(_GEN_26533); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26535 = 12'h3bb == _T_837 ? $signed(7'sh16) : $signed(_GEN_26534); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26536 = 12'h3bc == _T_837 ? $signed(7'sh17) : $signed(_GEN_26535); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26537 = 12'h3bd == _T_837 ? $signed(7'sh18) : $signed(_GEN_26536); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26538 = 12'h3be == _T_837 ? $signed(7'sh18) : $signed(_GEN_26537); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26539 = 12'h3bf == _T_837 ? $signed(7'sh19) : $signed(_GEN_26538); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26540 = 12'h3c0 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26539); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26541 = 12'h3c1 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26540); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26542 = 12'h3c2 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26541); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26543 = 12'h3c3 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26542); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26544 = 12'h3c4 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26543); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26545 = 12'h3c5 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26544); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26546 = 12'h3c6 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_26545); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26547 = 12'h3c7 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26546); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26548 = 12'h3c8 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26547); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26549 = 12'h3c9 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26548); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26550 = 12'h3ca == _T_837 ? $signed(7'sh1) : $signed(_GEN_26549); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26551 = 12'h3cb == _T_837 ? $signed(7'sh2) : $signed(_GEN_26550); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26552 = 12'h3cc == _T_837 ? $signed(7'sh3) : $signed(_GEN_26551); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26553 = 12'h3cd == _T_837 ? $signed(7'sh3) : $signed(_GEN_26552); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26554 = 12'h3ce == _T_837 ? $signed(7'sh4) : $signed(_GEN_26553); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26555 = 12'h3cf == _T_837 ? $signed(7'sh5) : $signed(_GEN_26554); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26556 = 12'h3d0 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26555); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26557 = 12'h3d1 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26556); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26558 = 12'h3d2 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26557); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26559 = 12'h3d3 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26558); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26560 = 12'h3d4 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26559); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26561 = 12'h3d5 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26560); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26562 = 12'h3d6 == _T_837 ? $signed(7'sha) : $signed(_GEN_26561); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26563 = 12'h3d7 == _T_837 ? $signed(7'sha) : $signed(_GEN_26562); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26564 = 12'h3d8 == _T_837 ? $signed(7'shb) : $signed(_GEN_26563); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26565 = 12'h3d9 == _T_837 ? $signed(7'shc) : $signed(_GEN_26564); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26566 = 12'h3da == _T_837 ? $signed(7'shc) : $signed(_GEN_26565); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26567 = 12'h3db == _T_837 ? $signed(7'shd) : $signed(_GEN_26566); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26568 = 12'h3dc == _T_837 ? $signed(7'she) : $signed(_GEN_26567); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26569 = 12'h3dd == _T_837 ? $signed(7'shf) : $signed(_GEN_26568); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26570 = 12'h3de == _T_837 ? $signed(7'shf) : $signed(_GEN_26569); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26571 = 12'h3df == _T_837 ? $signed(7'sh10) : $signed(_GEN_26570); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26572 = 12'h3e0 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26571); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26573 = 12'h3e1 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26572); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26574 = 12'h3e2 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26573); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26575 = 12'h3e3 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26574); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26576 = 12'h3e4 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26575); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26577 = 12'h3e5 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26576); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26578 = 12'h3e6 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26577); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26579 = 12'h3e7 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26578); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26580 = 12'h3e8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26579); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26581 = 12'h3e9 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26580); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26582 = 12'h3ea == _T_837 ? $signed(7'sh18) : $signed(_GEN_26581); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26583 = 12'h3eb == _T_837 ? $signed(7'sh18) : $signed(_GEN_26582); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26584 = 12'h3ec == _T_837 ? $signed(7'sh19) : $signed(_GEN_26583); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26585 = 12'h3ed == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26584); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26586 = 12'h3ee == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26585); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26587 = 12'h3ef == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26586); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26588 = 12'h3f0 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26587); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26589 = 12'h3f1 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26588); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26590 = 12'h3f2 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26589); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26591 = 12'h3f3 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26590); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26592 = 12'h3f4 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_26591); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26593 = 12'h3f5 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26592); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26594 = 12'h3f6 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26593); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26595 = 12'h3f7 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26594); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26596 = 12'h3f8 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26595); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26597 = 12'h3f9 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26596); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26598 = 12'h3fa == _T_837 ? $signed(7'sh3) : $signed(_GEN_26597); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26599 = 12'h3fb == _T_837 ? $signed(7'sh4) : $signed(_GEN_26598); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26600 = 12'h3fc == _T_837 ? $signed(7'sh5) : $signed(_GEN_26599); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26601 = 12'h3fd == _T_837 ? $signed(7'sh5) : $signed(_GEN_26600); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26602 = 12'h3fe == _T_837 ? $signed(7'sh6) : $signed(_GEN_26601); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26603 = 12'h3ff == _T_837 ? $signed(7'sh7) : $signed(_GEN_26602); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26604 = 12'h400 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26603); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26605 = 12'h401 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26604); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26606 = 12'h402 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26605); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26607 = 12'h403 == _T_837 ? $signed(7'sha) : $signed(_GEN_26606); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26608 = 12'h404 == _T_837 ? $signed(7'sha) : $signed(_GEN_26607); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26609 = 12'h405 == _T_837 ? $signed(7'shb) : $signed(_GEN_26608); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26610 = 12'h406 == _T_837 ? $signed(7'shc) : $signed(_GEN_26609); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26611 = 12'h407 == _T_837 ? $signed(7'shc) : $signed(_GEN_26610); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26612 = 12'h408 == _T_837 ? $signed(7'shd) : $signed(_GEN_26611); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26613 = 12'h409 == _T_837 ? $signed(7'she) : $signed(_GEN_26612); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26614 = 12'h40a == _T_837 ? $signed(7'shf) : $signed(_GEN_26613); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26615 = 12'h40b == _T_837 ? $signed(7'shf) : $signed(_GEN_26614); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26616 = 12'h40c == _T_837 ? $signed(7'sh10) : $signed(_GEN_26615); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26617 = 12'h40d == _T_837 ? $signed(7'sh11) : $signed(_GEN_26616); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26618 = 12'h40e == _T_837 ? $signed(7'sh11) : $signed(_GEN_26617); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26619 = 12'h40f == _T_837 ? $signed(7'sh12) : $signed(_GEN_26618); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26620 = 12'h410 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26619); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26621 = 12'h411 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26620); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26622 = 12'h412 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26621); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26623 = 12'h413 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26622); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26624 = 12'h414 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26623); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26625 = 12'h415 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26624); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26626 = 12'h416 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26625); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26627 = 12'h417 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26626); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26628 = 12'h418 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26627); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26629 = 12'h419 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26628); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26630 = 12'h41a == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26629); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26631 = 12'h41b == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26630); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26632 = 12'h41c == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26631); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26633 = 12'h41d == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26632); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26634 = 12'h41e == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26633); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26635 = 12'h41f == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26634); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26636 = 12'h420 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26635); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26637 = 12'h421 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26636); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26638 = 12'h422 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26637); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26639 = 12'h423 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26638); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26640 = 12'h424 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26639); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26641 = 12'h425 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26640); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26642 = 12'h426 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26641); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26643 = 12'h427 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26642); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26644 = 12'h428 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26643); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26645 = 12'h429 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26644); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26646 = 12'h42a == _T_837 ? $signed(7'sh5) : $signed(_GEN_26645); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26647 = 12'h42b == _T_837 ? $signed(7'sh6) : $signed(_GEN_26646); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26648 = 12'h42c == _T_837 ? $signed(7'sh7) : $signed(_GEN_26647); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26649 = 12'h42d == _T_837 ? $signed(7'sh8) : $signed(_GEN_26648); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26650 = 12'h42e == _T_837 ? $signed(7'sh8) : $signed(_GEN_26649); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26651 = 12'h42f == _T_837 ? $signed(7'sh9) : $signed(_GEN_26650); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26652 = 12'h430 == _T_837 ? $signed(7'sha) : $signed(_GEN_26651); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26653 = 12'h431 == _T_837 ? $signed(7'sha) : $signed(_GEN_26652); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26654 = 12'h432 == _T_837 ? $signed(7'shb) : $signed(_GEN_26653); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26655 = 12'h433 == _T_837 ? $signed(7'shc) : $signed(_GEN_26654); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26656 = 12'h434 == _T_837 ? $signed(7'shc) : $signed(_GEN_26655); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26657 = 12'h435 == _T_837 ? $signed(7'shd) : $signed(_GEN_26656); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26658 = 12'h436 == _T_837 ? $signed(7'she) : $signed(_GEN_26657); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26659 = 12'h437 == _T_837 ? $signed(7'shf) : $signed(_GEN_26658); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26660 = 12'h438 == _T_837 ? $signed(7'shf) : $signed(_GEN_26659); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26661 = 12'h439 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26660); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26662 = 12'h43a == _T_837 ? $signed(7'sh11) : $signed(_GEN_26661); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26663 = 12'h43b == _T_837 ? $signed(7'sh11) : $signed(_GEN_26662); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26664 = 12'h43c == _T_837 ? $signed(7'sh12) : $signed(_GEN_26663); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26665 = 12'h43d == _T_837 ? $signed(7'sh13) : $signed(_GEN_26664); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26666 = 12'h43e == _T_837 ? $signed(7'sh14) : $signed(_GEN_26665); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26667 = 12'h43f == _T_837 ? $signed(7'sh14) : $signed(_GEN_26666); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26668 = 12'h440 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26667); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26669 = 12'h441 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26668); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26670 = 12'h442 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26669); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26671 = 12'h443 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26670); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26672 = 12'h444 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26671); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26673 = 12'h445 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26672); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26674 = 12'h446 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26673); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26675 = 12'h447 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26674); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26676 = 12'h448 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26675); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26677 = 12'h449 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26676); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26678 = 12'h44a == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26677); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26679 = 12'h44b == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26678); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26680 = 12'h44c == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26679); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26681 = 12'h44d == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26680); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26682 = 12'h44e == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26681); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26683 = 12'h44f == _T_837 ? $signed(7'sh20) : $signed(_GEN_26682); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26684 = 12'h450 == _T_837 ? $signed(7'sh0) : $signed(_GEN_26683); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26685 = 12'h451 == _T_837 ? $signed(7'sh1) : $signed(_GEN_26684); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26686 = 12'h452 == _T_837 ? $signed(7'sh2) : $signed(_GEN_26685); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26687 = 12'h453 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26686); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26688 = 12'h454 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26687); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26689 = 12'h455 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26688); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26690 = 12'h456 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26689); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26691 = 12'h457 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26690); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26692 = 12'h458 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26691); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26693 = 12'h459 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26692); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26694 = 12'h45a == _T_837 ? $signed(7'sh8) : $signed(_GEN_26693); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26695 = 12'h45b == _T_837 ? $signed(7'sh8) : $signed(_GEN_26694); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26696 = 12'h45c == _T_837 ? $signed(7'sh9) : $signed(_GEN_26695); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26697 = 12'h45d == _T_837 ? $signed(7'sha) : $signed(_GEN_26696); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26698 = 12'h45e == _T_837 ? $signed(7'sha) : $signed(_GEN_26697); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26699 = 12'h45f == _T_837 ? $signed(7'shb) : $signed(_GEN_26698); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26700 = 12'h460 == _T_837 ? $signed(7'shc) : $signed(_GEN_26699); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26701 = 12'h461 == _T_837 ? $signed(7'shc) : $signed(_GEN_26700); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26702 = 12'h462 == _T_837 ? $signed(7'shd) : $signed(_GEN_26701); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26703 = 12'h463 == _T_837 ? $signed(7'she) : $signed(_GEN_26702); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26704 = 12'h464 == _T_837 ? $signed(7'shf) : $signed(_GEN_26703); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26705 = 12'h465 == _T_837 ? $signed(7'shf) : $signed(_GEN_26704); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26706 = 12'h466 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26705); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26707 = 12'h467 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26706); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26708 = 12'h468 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26707); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26709 = 12'h469 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26708); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26710 = 12'h46a == _T_837 ? $signed(7'sh13) : $signed(_GEN_26709); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26711 = 12'h46b == _T_837 ? $signed(7'sh14) : $signed(_GEN_26710); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26712 = 12'h46c == _T_837 ? $signed(7'sh14) : $signed(_GEN_26711); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26713 = 12'h46d == _T_837 ? $signed(7'sh15) : $signed(_GEN_26712); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26714 = 12'h46e == _T_837 ? $signed(7'sh16) : $signed(_GEN_26713); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26715 = 12'h46f == _T_837 ? $signed(7'sh16) : $signed(_GEN_26714); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26716 = 12'h470 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26715); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26717 = 12'h471 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26716); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26718 = 12'h472 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26717); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26719 = 12'h473 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26718); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26720 = 12'h474 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26719); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26721 = 12'h475 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26720); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26722 = 12'h476 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26721); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26723 = 12'h477 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26722); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26724 = 12'h478 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26723); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26725 = 12'h479 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26724); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26726 = 12'h47a == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26725); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26727 = 12'h47b == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26726); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26728 = 12'h47c == _T_837 ? $signed(7'sh20) : $signed(_GEN_26727); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26729 = 12'h47d == _T_837 ? $signed(7'sh20) : $signed(_GEN_26728); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26730 = 12'h47e == _T_837 ? $signed(7'sh1) : $signed(_GEN_26729); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26731 = 12'h47f == _T_837 ? $signed(7'sh2) : $signed(_GEN_26730); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26732 = 12'h480 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26731); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26733 = 12'h481 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26732); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26734 = 12'h482 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26733); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26735 = 12'h483 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26734); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26736 = 12'h484 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26735); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26737 = 12'h485 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26736); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26738 = 12'h486 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26737); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26739 = 12'h487 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26738); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26740 = 12'h488 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26739); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26741 = 12'h489 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26740); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26742 = 12'h48a == _T_837 ? $signed(7'sha) : $signed(_GEN_26741); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26743 = 12'h48b == _T_837 ? $signed(7'sha) : $signed(_GEN_26742); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26744 = 12'h48c == _T_837 ? $signed(7'shb) : $signed(_GEN_26743); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26745 = 12'h48d == _T_837 ? $signed(7'shc) : $signed(_GEN_26744); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26746 = 12'h48e == _T_837 ? $signed(7'shc) : $signed(_GEN_26745); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26747 = 12'h48f == _T_837 ? $signed(7'shd) : $signed(_GEN_26746); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26748 = 12'h490 == _T_837 ? $signed(7'she) : $signed(_GEN_26747); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26749 = 12'h491 == _T_837 ? $signed(7'shf) : $signed(_GEN_26748); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26750 = 12'h492 == _T_837 ? $signed(7'shf) : $signed(_GEN_26749); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26751 = 12'h493 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26750); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26752 = 12'h494 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26751); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26753 = 12'h495 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26752); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26754 = 12'h496 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26753); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26755 = 12'h497 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26754); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26756 = 12'h498 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26755); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26757 = 12'h499 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26756); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26758 = 12'h49a == _T_837 ? $signed(7'sh15) : $signed(_GEN_26757); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26759 = 12'h49b == _T_837 ? $signed(7'sh16) : $signed(_GEN_26758); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26760 = 12'h49c == _T_837 ? $signed(7'sh16) : $signed(_GEN_26759); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26761 = 12'h49d == _T_837 ? $signed(7'sh17) : $signed(_GEN_26760); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26762 = 12'h49e == _T_837 ? $signed(7'sh18) : $signed(_GEN_26761); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26763 = 12'h49f == _T_837 ? $signed(7'sh18) : $signed(_GEN_26762); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26764 = 12'h4a0 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26763); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26765 = 12'h4a1 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26764); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26766 = 12'h4a2 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26765); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26767 = 12'h4a3 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26766); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26768 = 12'h4a4 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26767); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26769 = 12'h4a5 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26768); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26770 = 12'h4a6 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26769); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26771 = 12'h4a7 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26770); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26772 = 12'h4a8 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26771); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26773 = 12'h4a9 == _T_837 ? $signed(7'sh20) : $signed(_GEN_26772); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26774 = 12'h4aa == _T_837 ? $signed(7'sh20) : $signed(_GEN_26773); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26775 = 12'h4ab == _T_837 ? $signed(7'sh21) : $signed(_GEN_26774); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26776 = 12'h4ac == _T_837 ? $signed(7'sh2) : $signed(_GEN_26775); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26777 = 12'h4ad == _T_837 ? $signed(7'sh3) : $signed(_GEN_26776); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26778 = 12'h4ae == _T_837 ? $signed(7'sh3) : $signed(_GEN_26777); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26779 = 12'h4af == _T_837 ? $signed(7'sh4) : $signed(_GEN_26778); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26780 = 12'h4b0 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26779); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26781 = 12'h4b1 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26780); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26782 = 12'h4b2 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26781); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26783 = 12'h4b3 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26782); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26784 = 12'h4b4 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26783); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26785 = 12'h4b5 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26784); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26786 = 12'h4b6 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26785); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26787 = 12'h4b7 == _T_837 ? $signed(7'sha) : $signed(_GEN_26786); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26788 = 12'h4b8 == _T_837 ? $signed(7'sha) : $signed(_GEN_26787); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26789 = 12'h4b9 == _T_837 ? $signed(7'shb) : $signed(_GEN_26788); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26790 = 12'h4ba == _T_837 ? $signed(7'shc) : $signed(_GEN_26789); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26791 = 12'h4bb == _T_837 ? $signed(7'shc) : $signed(_GEN_26790); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26792 = 12'h4bc == _T_837 ? $signed(7'shd) : $signed(_GEN_26791); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26793 = 12'h4bd == _T_837 ? $signed(7'she) : $signed(_GEN_26792); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26794 = 12'h4be == _T_837 ? $signed(7'shf) : $signed(_GEN_26793); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26795 = 12'h4bf == _T_837 ? $signed(7'shf) : $signed(_GEN_26794); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26796 = 12'h4c0 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26795); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26797 = 12'h4c1 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26796); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26798 = 12'h4c2 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26797); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26799 = 12'h4c3 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26798); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26800 = 12'h4c4 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26799); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26801 = 12'h4c5 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26800); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26802 = 12'h4c6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26801); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26803 = 12'h4c7 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26802); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26804 = 12'h4c8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26803); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26805 = 12'h4c9 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26804); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26806 = 12'h4ca == _T_837 ? $signed(7'sh17) : $signed(_GEN_26805); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26807 = 12'h4cb == _T_837 ? $signed(7'sh18) : $signed(_GEN_26806); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26808 = 12'h4cc == _T_837 ? $signed(7'sh18) : $signed(_GEN_26807); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26809 = 12'h4cd == _T_837 ? $signed(7'sh19) : $signed(_GEN_26808); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26810 = 12'h4ce == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26809); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26811 = 12'h4cf == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26810); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26812 = 12'h4d0 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26811); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26813 = 12'h4d1 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26812); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26814 = 12'h4d2 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26813); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26815 = 12'h4d3 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26814); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26816 = 12'h4d4 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26815); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26817 = 12'h4d5 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26816); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26818 = 12'h4d6 == _T_837 ? $signed(7'sh20) : $signed(_GEN_26817); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26819 = 12'h4d7 == _T_837 ? $signed(7'sh20) : $signed(_GEN_26818); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26820 = 12'h4d8 == _T_837 ? $signed(7'sh21) : $signed(_GEN_26819); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26821 = 12'h4d9 == _T_837 ? $signed(7'sh22) : $signed(_GEN_26820); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26822 = 12'h4da == _T_837 ? $signed(7'sh3) : $signed(_GEN_26821); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26823 = 12'h4db == _T_837 ? $signed(7'sh3) : $signed(_GEN_26822); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26824 = 12'h4dc == _T_837 ? $signed(7'sh4) : $signed(_GEN_26823); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26825 = 12'h4dd == _T_837 ? $signed(7'sh5) : $signed(_GEN_26824); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26826 = 12'h4de == _T_837 ? $signed(7'sh5) : $signed(_GEN_26825); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26827 = 12'h4df == _T_837 ? $signed(7'sh6) : $signed(_GEN_26826); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26828 = 12'h4e0 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26827); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26829 = 12'h4e1 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26828); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26830 = 12'h4e2 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26829); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26831 = 12'h4e3 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26830); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26832 = 12'h4e4 == _T_837 ? $signed(7'sha) : $signed(_GEN_26831); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26833 = 12'h4e5 == _T_837 ? $signed(7'sha) : $signed(_GEN_26832); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26834 = 12'h4e6 == _T_837 ? $signed(7'shb) : $signed(_GEN_26833); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26835 = 12'h4e7 == _T_837 ? $signed(7'shc) : $signed(_GEN_26834); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26836 = 12'h4e8 == _T_837 ? $signed(7'shc) : $signed(_GEN_26835); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26837 = 12'h4e9 == _T_837 ? $signed(7'shd) : $signed(_GEN_26836); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26838 = 12'h4ea == _T_837 ? $signed(7'she) : $signed(_GEN_26837); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26839 = 12'h4eb == _T_837 ? $signed(7'shf) : $signed(_GEN_26838); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26840 = 12'h4ec == _T_837 ? $signed(7'shf) : $signed(_GEN_26839); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26841 = 12'h4ed == _T_837 ? $signed(7'sh10) : $signed(_GEN_26840); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26842 = 12'h4ee == _T_837 ? $signed(7'sh11) : $signed(_GEN_26841); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26843 = 12'h4ef == _T_837 ? $signed(7'sh11) : $signed(_GEN_26842); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26844 = 12'h4f0 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26843); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26845 = 12'h4f1 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26844); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26846 = 12'h4f2 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26845); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26847 = 12'h4f3 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26846); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26848 = 12'h4f4 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26847); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26849 = 12'h4f5 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26848); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26850 = 12'h4f6 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26849); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26851 = 12'h4f7 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26850); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26852 = 12'h4f8 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26851); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26853 = 12'h4f9 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26852); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26854 = 12'h4fa == _T_837 ? $signed(7'sh19) : $signed(_GEN_26853); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26855 = 12'h4fb == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26854); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26856 = 12'h4fc == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26855); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26857 = 12'h4fd == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26856); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26858 = 12'h4fe == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26857); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26859 = 12'h4ff == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26858); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26860 = 12'h500 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26859); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26861 = 12'h501 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26860); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26862 = 12'h502 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26861); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26863 = 12'h503 == _T_837 ? $signed(7'sh20) : $signed(_GEN_26862); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26864 = 12'h504 == _T_837 ? $signed(7'sh20) : $signed(_GEN_26863); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26865 = 12'h505 == _T_837 ? $signed(7'sh21) : $signed(_GEN_26864); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26866 = 12'h506 == _T_837 ? $signed(7'sh22) : $signed(_GEN_26865); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26867 = 12'h507 == _T_837 ? $signed(7'sh22) : $signed(_GEN_26866); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26868 = 12'h508 == _T_837 ? $signed(7'sh3) : $signed(_GEN_26867); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26869 = 12'h509 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26868); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26870 = 12'h50a == _T_837 ? $signed(7'sh5) : $signed(_GEN_26869); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26871 = 12'h50b == _T_837 ? $signed(7'sh5) : $signed(_GEN_26870); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26872 = 12'h50c == _T_837 ? $signed(7'sh6) : $signed(_GEN_26871); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26873 = 12'h50d == _T_837 ? $signed(7'sh7) : $signed(_GEN_26872); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26874 = 12'h50e == _T_837 ? $signed(7'sh8) : $signed(_GEN_26873); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26875 = 12'h50f == _T_837 ? $signed(7'sh8) : $signed(_GEN_26874); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26876 = 12'h510 == _T_837 ? $signed(7'sh9) : $signed(_GEN_26875); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26877 = 12'h511 == _T_837 ? $signed(7'sha) : $signed(_GEN_26876); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26878 = 12'h512 == _T_837 ? $signed(7'sha) : $signed(_GEN_26877); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26879 = 12'h513 == _T_837 ? $signed(7'shb) : $signed(_GEN_26878); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26880 = 12'h514 == _T_837 ? $signed(7'shc) : $signed(_GEN_26879); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26881 = 12'h515 == _T_837 ? $signed(7'shc) : $signed(_GEN_26880); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26882 = 12'h516 == _T_837 ? $signed(7'shd) : $signed(_GEN_26881); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26883 = 12'h517 == _T_837 ? $signed(7'she) : $signed(_GEN_26882); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26884 = 12'h518 == _T_837 ? $signed(7'shf) : $signed(_GEN_26883); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26885 = 12'h519 == _T_837 ? $signed(7'shf) : $signed(_GEN_26884); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26886 = 12'h51a == _T_837 ? $signed(7'sh10) : $signed(_GEN_26885); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26887 = 12'h51b == _T_837 ? $signed(7'sh11) : $signed(_GEN_26886); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26888 = 12'h51c == _T_837 ? $signed(7'sh11) : $signed(_GEN_26887); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26889 = 12'h51d == _T_837 ? $signed(7'sh12) : $signed(_GEN_26888); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26890 = 12'h51e == _T_837 ? $signed(7'sh13) : $signed(_GEN_26889); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26891 = 12'h51f == _T_837 ? $signed(7'sh14) : $signed(_GEN_26890); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26892 = 12'h520 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26891); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26893 = 12'h521 == _T_837 ? $signed(7'sh15) : $signed(_GEN_26892); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26894 = 12'h522 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26893); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26895 = 12'h523 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26894); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26896 = 12'h524 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26895); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26897 = 12'h525 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26896); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26898 = 12'h526 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26897); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26899 = 12'h527 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26898); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26900 = 12'h528 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26899); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26901 = 12'h529 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26900); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26902 = 12'h52a == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26901); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26903 = 12'h52b == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26902); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26904 = 12'h52c == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26903); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26905 = 12'h52d == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26904); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26906 = 12'h52e == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26905); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26907 = 12'h52f == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26906); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26908 = 12'h530 == _T_837 ? $signed(7'sh20) : $signed(_GEN_26907); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26909 = 12'h531 == _T_837 ? $signed(7'sh20) : $signed(_GEN_26908); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26910 = 12'h532 == _T_837 ? $signed(7'sh21) : $signed(_GEN_26909); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26911 = 12'h533 == _T_837 ? $signed(7'sh22) : $signed(_GEN_26910); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26912 = 12'h534 == _T_837 ? $signed(7'sh22) : $signed(_GEN_26911); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26913 = 12'h535 == _T_837 ? $signed(7'sh23) : $signed(_GEN_26912); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26914 = 12'h536 == _T_837 ? $signed(7'sh4) : $signed(_GEN_26913); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26915 = 12'h537 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26914); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26916 = 12'h538 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26915); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26917 = 12'h539 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26916); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26918 = 12'h53a == _T_837 ? $signed(7'sh7) : $signed(_GEN_26917); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26919 = 12'h53b == _T_837 ? $signed(7'sh8) : $signed(_GEN_26918); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26920 = 12'h53c == _T_837 ? $signed(7'sh8) : $signed(_GEN_26919); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26921 = 12'h53d == _T_837 ? $signed(7'sh9) : $signed(_GEN_26920); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26922 = 12'h53e == _T_837 ? $signed(7'sha) : $signed(_GEN_26921); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26923 = 12'h53f == _T_837 ? $signed(7'sha) : $signed(_GEN_26922); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26924 = 12'h540 == _T_837 ? $signed(7'shb) : $signed(_GEN_26923); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26925 = 12'h541 == _T_837 ? $signed(7'shc) : $signed(_GEN_26924); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26926 = 12'h542 == _T_837 ? $signed(7'shc) : $signed(_GEN_26925); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26927 = 12'h543 == _T_837 ? $signed(7'shd) : $signed(_GEN_26926); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26928 = 12'h544 == _T_837 ? $signed(7'she) : $signed(_GEN_26927); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26929 = 12'h545 == _T_837 ? $signed(7'shf) : $signed(_GEN_26928); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26930 = 12'h546 == _T_837 ? $signed(7'shf) : $signed(_GEN_26929); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26931 = 12'h547 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26930); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26932 = 12'h548 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26931); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26933 = 12'h549 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26932); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26934 = 12'h54a == _T_837 ? $signed(7'sh12) : $signed(_GEN_26933); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26935 = 12'h54b == _T_837 ? $signed(7'sh13) : $signed(_GEN_26934); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26936 = 12'h54c == _T_837 ? $signed(7'sh14) : $signed(_GEN_26935); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26937 = 12'h54d == _T_837 ? $signed(7'sh14) : $signed(_GEN_26936); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26938 = 12'h54e == _T_837 ? $signed(7'sh15) : $signed(_GEN_26937); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26939 = 12'h54f == _T_837 ? $signed(7'sh16) : $signed(_GEN_26938); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26940 = 12'h550 == _T_837 ? $signed(7'sh16) : $signed(_GEN_26939); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26941 = 12'h551 == _T_837 ? $signed(7'sh17) : $signed(_GEN_26940); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26942 = 12'h552 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26941); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26943 = 12'h553 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26942); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26944 = 12'h554 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26943); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26945 = 12'h555 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26944); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26946 = 12'h556 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26945); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26947 = 12'h557 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26946); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26948 = 12'h558 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26947); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26949 = 12'h559 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26948); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26950 = 12'h55a == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26949); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26951 = 12'h55b == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26950); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26952 = 12'h55c == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26951); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26953 = 12'h55d == _T_837 ? $signed(7'sh20) : $signed(_GEN_26952); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26954 = 12'h55e == _T_837 ? $signed(7'sh20) : $signed(_GEN_26953); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26955 = 12'h55f == _T_837 ? $signed(7'sh21) : $signed(_GEN_26954); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26956 = 12'h560 == _T_837 ? $signed(7'sh22) : $signed(_GEN_26955); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26957 = 12'h561 == _T_837 ? $signed(7'sh22) : $signed(_GEN_26956); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26958 = 12'h562 == _T_837 ? $signed(7'sh23) : $signed(_GEN_26957); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26959 = 12'h563 == _T_837 ? $signed(7'sh24) : $signed(_GEN_26958); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26960 = 12'h564 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26959); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26961 = 12'h565 == _T_837 ? $signed(7'sh5) : $signed(_GEN_26960); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26962 = 12'h566 == _T_837 ? $signed(7'sh6) : $signed(_GEN_26961); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26963 = 12'h567 == _T_837 ? $signed(7'sh7) : $signed(_GEN_26962); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26964 = 12'h568 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26963); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26965 = 12'h569 == _T_837 ? $signed(7'sh8) : $signed(_GEN_26964); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26966 = 12'h56a == _T_837 ? $signed(7'sh9) : $signed(_GEN_26965); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26967 = 12'h56b == _T_837 ? $signed(7'sha) : $signed(_GEN_26966); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26968 = 12'h56c == _T_837 ? $signed(7'sha) : $signed(_GEN_26967); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26969 = 12'h56d == _T_837 ? $signed(7'shb) : $signed(_GEN_26968); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26970 = 12'h56e == _T_837 ? $signed(7'shc) : $signed(_GEN_26969); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26971 = 12'h56f == _T_837 ? $signed(7'shc) : $signed(_GEN_26970); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26972 = 12'h570 == _T_837 ? $signed(7'shd) : $signed(_GEN_26971); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26973 = 12'h571 == _T_837 ? $signed(7'she) : $signed(_GEN_26972); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26974 = 12'h572 == _T_837 ? $signed(7'shf) : $signed(_GEN_26973); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26975 = 12'h573 == _T_837 ? $signed(7'shf) : $signed(_GEN_26974); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26976 = 12'h574 == _T_837 ? $signed(7'sh10) : $signed(_GEN_26975); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26977 = 12'h575 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26976); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26978 = 12'h576 == _T_837 ? $signed(7'sh11) : $signed(_GEN_26977); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26979 = 12'h577 == _T_837 ? $signed(7'sh12) : $signed(_GEN_26978); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26980 = 12'h578 == _T_837 ? $signed(7'sh13) : $signed(_GEN_26979); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26981 = 12'h579 == _T_837 ? $signed(7'sh14) : $signed(_GEN_26980); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26982 = 12'h57a == _T_837 ? $signed(7'sh14) : $signed(_GEN_26981); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26983 = 12'h57b == _T_837 ? $signed(7'sh15) : $signed(_GEN_26982); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26984 = 12'h57c == _T_837 ? $signed(7'sh16) : $signed(_GEN_26983); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26985 = 12'h57d == _T_837 ? $signed(7'sh16) : $signed(_GEN_26984); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26986 = 12'h57e == _T_837 ? $signed(7'sh17) : $signed(_GEN_26985); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26987 = 12'h57f == _T_837 ? $signed(7'sh18) : $signed(_GEN_26986); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26988 = 12'h580 == _T_837 ? $signed(7'sh18) : $signed(_GEN_26987); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26989 = 12'h581 == _T_837 ? $signed(7'sh19) : $signed(_GEN_26988); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26990 = 12'h582 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_26989); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26991 = 12'h583 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26990); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26992 = 12'h584 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_26991); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26993 = 12'h585 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_26992); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26994 = 12'h586 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26993); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26995 = 12'h587 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_26994); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26996 = 12'h588 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_26995); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26997 = 12'h589 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_26996); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26998 = 12'h58a == _T_837 ? $signed(7'sh20) : $signed(_GEN_26997); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_26999 = 12'h58b == _T_837 ? $signed(7'sh20) : $signed(_GEN_26998); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27000 = 12'h58c == _T_837 ? $signed(7'sh21) : $signed(_GEN_26999); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27001 = 12'h58d == _T_837 ? $signed(7'sh22) : $signed(_GEN_27000); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27002 = 12'h58e == _T_837 ? $signed(7'sh22) : $signed(_GEN_27001); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27003 = 12'h58f == _T_837 ? $signed(7'sh23) : $signed(_GEN_27002); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27004 = 12'h590 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27003); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27005 = 12'h591 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27004); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27006 = 12'h592 == _T_837 ? $signed(7'sh5) : $signed(_GEN_27005); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27007 = 12'h593 == _T_837 ? $signed(7'sh6) : $signed(_GEN_27006); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27008 = 12'h594 == _T_837 ? $signed(7'sh7) : $signed(_GEN_27007); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27009 = 12'h595 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27008); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27010 = 12'h596 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27009); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27011 = 12'h597 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27010); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27012 = 12'h598 == _T_837 ? $signed(7'sha) : $signed(_GEN_27011); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27013 = 12'h599 == _T_837 ? $signed(7'sha) : $signed(_GEN_27012); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27014 = 12'h59a == _T_837 ? $signed(7'shb) : $signed(_GEN_27013); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27015 = 12'h59b == _T_837 ? $signed(7'shc) : $signed(_GEN_27014); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27016 = 12'h59c == _T_837 ? $signed(7'shc) : $signed(_GEN_27015); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27017 = 12'h59d == _T_837 ? $signed(7'shd) : $signed(_GEN_27016); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27018 = 12'h59e == _T_837 ? $signed(7'she) : $signed(_GEN_27017); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27019 = 12'h59f == _T_837 ? $signed(7'shf) : $signed(_GEN_27018); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27020 = 12'h5a0 == _T_837 ? $signed(7'shf) : $signed(_GEN_27019); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27021 = 12'h5a1 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27020); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27022 = 12'h5a2 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27021); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27023 = 12'h5a3 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27022); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27024 = 12'h5a4 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27023); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27025 = 12'h5a5 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27024); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27026 = 12'h5a6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27025); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27027 = 12'h5a7 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27026); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27028 = 12'h5a8 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27027); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27029 = 12'h5a9 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27028); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27030 = 12'h5aa == _T_837 ? $signed(7'sh16) : $signed(_GEN_27029); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27031 = 12'h5ab == _T_837 ? $signed(7'sh17) : $signed(_GEN_27030); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27032 = 12'h5ac == _T_837 ? $signed(7'sh18) : $signed(_GEN_27031); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27033 = 12'h5ad == _T_837 ? $signed(7'sh18) : $signed(_GEN_27032); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27034 = 12'h5ae == _T_837 ? $signed(7'sh19) : $signed(_GEN_27033); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27035 = 12'h5af == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27034); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27036 = 12'h5b0 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27035); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27037 = 12'h5b1 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27036); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27038 = 12'h5b2 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27037); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27039 = 12'h5b3 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27038); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27040 = 12'h5b4 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27039); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27041 = 12'h5b5 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27040); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27042 = 12'h5b6 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27041); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27043 = 12'h5b7 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27042); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27044 = 12'h5b8 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27043); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27045 = 12'h5b9 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27044); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27046 = 12'h5ba == _T_837 ? $signed(7'sh22) : $signed(_GEN_27045); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27047 = 12'h5bb == _T_837 ? $signed(7'sh22) : $signed(_GEN_27046); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27048 = 12'h5bc == _T_837 ? $signed(7'sh23) : $signed(_GEN_27047); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27049 = 12'h5bd == _T_837 ? $signed(7'sh24) : $signed(_GEN_27048); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27050 = 12'h5be == _T_837 ? $signed(7'sh25) : $signed(_GEN_27049); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27051 = 12'h5bf == _T_837 ? $signed(7'sh25) : $signed(_GEN_27050); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27052 = 12'h5c0 == _T_837 ? $signed(7'sh6) : $signed(_GEN_27051); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27053 = 12'h5c1 == _T_837 ? $signed(7'sh7) : $signed(_GEN_27052); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27054 = 12'h5c2 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27053); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27055 = 12'h5c3 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27054); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27056 = 12'h5c4 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27055); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27057 = 12'h5c5 == _T_837 ? $signed(7'sha) : $signed(_GEN_27056); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27058 = 12'h5c6 == _T_837 ? $signed(7'sha) : $signed(_GEN_27057); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27059 = 12'h5c7 == _T_837 ? $signed(7'shb) : $signed(_GEN_27058); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27060 = 12'h5c8 == _T_837 ? $signed(7'shc) : $signed(_GEN_27059); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27061 = 12'h5c9 == _T_837 ? $signed(7'shc) : $signed(_GEN_27060); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27062 = 12'h5ca == _T_837 ? $signed(7'shd) : $signed(_GEN_27061); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27063 = 12'h5cb == _T_837 ? $signed(7'she) : $signed(_GEN_27062); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27064 = 12'h5cc == _T_837 ? $signed(7'shf) : $signed(_GEN_27063); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27065 = 12'h5cd == _T_837 ? $signed(7'shf) : $signed(_GEN_27064); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27066 = 12'h5ce == _T_837 ? $signed(7'sh10) : $signed(_GEN_27065); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27067 = 12'h5cf == _T_837 ? $signed(7'sh11) : $signed(_GEN_27066); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27068 = 12'h5d0 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27067); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27069 = 12'h5d1 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27068); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27070 = 12'h5d2 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27069); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27071 = 12'h5d3 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27070); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27072 = 12'h5d4 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27071); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27073 = 12'h5d5 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27072); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27074 = 12'h5d6 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27073); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27075 = 12'h5d7 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27074); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27076 = 12'h5d8 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27075); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27077 = 12'h5d9 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27076); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27078 = 12'h5da == _T_837 ? $signed(7'sh18) : $signed(_GEN_27077); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27079 = 12'h5db == _T_837 ? $signed(7'sh19) : $signed(_GEN_27078); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27080 = 12'h5dc == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27079); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27081 = 12'h5dd == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27080); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27082 = 12'h5de == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27081); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27083 = 12'h5df == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27082); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27084 = 12'h5e0 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27083); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27085 = 12'h5e1 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27084); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27086 = 12'h5e2 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27085); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27087 = 12'h5e3 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27086); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27088 = 12'h5e4 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27087); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27089 = 12'h5e5 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27088); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27090 = 12'h5e6 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27089); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27091 = 12'h5e7 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27090); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27092 = 12'h5e8 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27091); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27093 = 12'h5e9 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27092); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27094 = 12'h5ea == _T_837 ? $signed(7'sh24) : $signed(_GEN_27093); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27095 = 12'h5eb == _T_837 ? $signed(7'sh25) : $signed(_GEN_27094); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27096 = 12'h5ec == _T_837 ? $signed(7'sh25) : $signed(_GEN_27095); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27097 = 12'h5ed == _T_837 ? $signed(7'sh26) : $signed(_GEN_27096); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27098 = 12'h5ee == _T_837 ? $signed(7'sh7) : $signed(_GEN_27097); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27099 = 12'h5ef == _T_837 ? $signed(7'sh8) : $signed(_GEN_27098); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27100 = 12'h5f0 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27099); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27101 = 12'h5f1 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27100); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27102 = 12'h5f2 == _T_837 ? $signed(7'sha) : $signed(_GEN_27101); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27103 = 12'h5f3 == _T_837 ? $signed(7'sha) : $signed(_GEN_27102); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27104 = 12'h5f4 == _T_837 ? $signed(7'shb) : $signed(_GEN_27103); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27105 = 12'h5f5 == _T_837 ? $signed(7'shc) : $signed(_GEN_27104); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27106 = 12'h5f6 == _T_837 ? $signed(7'shc) : $signed(_GEN_27105); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27107 = 12'h5f7 == _T_837 ? $signed(7'shd) : $signed(_GEN_27106); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27108 = 12'h5f8 == _T_837 ? $signed(7'she) : $signed(_GEN_27107); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27109 = 12'h5f9 == _T_837 ? $signed(7'shf) : $signed(_GEN_27108); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27110 = 12'h5fa == _T_837 ? $signed(7'shf) : $signed(_GEN_27109); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27111 = 12'h5fb == _T_837 ? $signed(7'sh10) : $signed(_GEN_27110); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27112 = 12'h5fc == _T_837 ? $signed(7'sh11) : $signed(_GEN_27111); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27113 = 12'h5fd == _T_837 ? $signed(7'sh11) : $signed(_GEN_27112); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27114 = 12'h5fe == _T_837 ? $signed(7'sh12) : $signed(_GEN_27113); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27115 = 12'h5ff == _T_837 ? $signed(7'sh13) : $signed(_GEN_27114); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27116 = 12'h600 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27115); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27117 = 12'h601 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27116); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27118 = 12'h602 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27117); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27119 = 12'h603 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27118); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27120 = 12'h604 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27119); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27121 = 12'h605 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27120); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27122 = 12'h606 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27121); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27123 = 12'h607 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27122); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27124 = 12'h608 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27123); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27125 = 12'h609 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27124); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27126 = 12'h60a == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27125); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27127 = 12'h60b == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27126); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27128 = 12'h60c == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27127); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27129 = 12'h60d == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27128); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27130 = 12'h60e == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27129); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27131 = 12'h60f == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27130); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27132 = 12'h610 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27131); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27133 = 12'h611 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27132); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27134 = 12'h612 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27133); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27135 = 12'h613 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27134); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27136 = 12'h614 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27135); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27137 = 12'h615 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27136); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27138 = 12'h616 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27137); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27139 = 12'h617 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27138); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27140 = 12'h618 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27139); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27141 = 12'h619 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27140); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27142 = 12'h61a == _T_837 ? $signed(7'sh26) : $signed(_GEN_27141); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27143 = 12'h61b == _T_837 ? $signed(7'sh27) : $signed(_GEN_27142); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27144 = 12'h61c == _T_837 ? $signed(7'sh8) : $signed(_GEN_27143); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27145 = 12'h61d == _T_837 ? $signed(7'sh8) : $signed(_GEN_27144); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27146 = 12'h61e == _T_837 ? $signed(7'sh9) : $signed(_GEN_27145); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27147 = 12'h61f == _T_837 ? $signed(7'sha) : $signed(_GEN_27146); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27148 = 12'h620 == _T_837 ? $signed(7'sha) : $signed(_GEN_27147); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27149 = 12'h621 == _T_837 ? $signed(7'shb) : $signed(_GEN_27148); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27150 = 12'h622 == _T_837 ? $signed(7'shc) : $signed(_GEN_27149); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27151 = 12'h623 == _T_837 ? $signed(7'shc) : $signed(_GEN_27150); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27152 = 12'h624 == _T_837 ? $signed(7'shd) : $signed(_GEN_27151); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27153 = 12'h625 == _T_837 ? $signed(7'she) : $signed(_GEN_27152); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27154 = 12'h626 == _T_837 ? $signed(7'shf) : $signed(_GEN_27153); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27155 = 12'h627 == _T_837 ? $signed(7'shf) : $signed(_GEN_27154); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27156 = 12'h628 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27155); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27157 = 12'h629 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27156); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27158 = 12'h62a == _T_837 ? $signed(7'sh11) : $signed(_GEN_27157); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27159 = 12'h62b == _T_837 ? $signed(7'sh12) : $signed(_GEN_27158); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27160 = 12'h62c == _T_837 ? $signed(7'sh13) : $signed(_GEN_27159); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27161 = 12'h62d == _T_837 ? $signed(7'sh14) : $signed(_GEN_27160); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27162 = 12'h62e == _T_837 ? $signed(7'sh14) : $signed(_GEN_27161); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27163 = 12'h62f == _T_837 ? $signed(7'sh15) : $signed(_GEN_27162); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27164 = 12'h630 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27163); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27165 = 12'h631 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27164); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27166 = 12'h632 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27165); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27167 = 12'h633 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27166); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27168 = 12'h634 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27167); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27169 = 12'h635 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27168); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27170 = 12'h636 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27169); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27171 = 12'h637 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27170); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27172 = 12'h638 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27171); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27173 = 12'h639 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27172); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27174 = 12'h63a == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27173); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27175 = 12'h63b == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27174); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27176 = 12'h63c == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27175); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27177 = 12'h63d == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27176); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27178 = 12'h63e == _T_837 ? $signed(7'sh20) : $signed(_GEN_27177); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27179 = 12'h63f == _T_837 ? $signed(7'sh20) : $signed(_GEN_27178); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27180 = 12'h640 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27179); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27181 = 12'h641 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27180); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27182 = 12'h642 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27181); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27183 = 12'h643 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27182); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27184 = 12'h644 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27183); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27185 = 12'h645 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27184); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27186 = 12'h646 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27185); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27187 = 12'h647 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27186); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27188 = 12'h648 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27187); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27189 = 12'h649 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27188); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27190 = 12'h64a == _T_837 ? $signed(7'sh8) : $signed(_GEN_27189); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27191 = 12'h64b == _T_837 ? $signed(7'sh9) : $signed(_GEN_27190); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27192 = 12'h64c == _T_837 ? $signed(7'sha) : $signed(_GEN_27191); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27193 = 12'h64d == _T_837 ? $signed(7'sha) : $signed(_GEN_27192); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27194 = 12'h64e == _T_837 ? $signed(7'shb) : $signed(_GEN_27193); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27195 = 12'h64f == _T_837 ? $signed(7'shc) : $signed(_GEN_27194); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27196 = 12'h650 == _T_837 ? $signed(7'shc) : $signed(_GEN_27195); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27197 = 12'h651 == _T_837 ? $signed(7'shd) : $signed(_GEN_27196); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27198 = 12'h652 == _T_837 ? $signed(7'she) : $signed(_GEN_27197); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27199 = 12'h653 == _T_837 ? $signed(7'shf) : $signed(_GEN_27198); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27200 = 12'h654 == _T_837 ? $signed(7'shf) : $signed(_GEN_27199); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27201 = 12'h655 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27200); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27202 = 12'h656 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27201); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27203 = 12'h657 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27202); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27204 = 12'h658 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27203); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27205 = 12'h659 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27204); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27206 = 12'h65a == _T_837 ? $signed(7'sh14) : $signed(_GEN_27205); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27207 = 12'h65b == _T_837 ? $signed(7'sh14) : $signed(_GEN_27206); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27208 = 12'h65c == _T_837 ? $signed(7'sh15) : $signed(_GEN_27207); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27209 = 12'h65d == _T_837 ? $signed(7'sh16) : $signed(_GEN_27208); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27210 = 12'h65e == _T_837 ? $signed(7'sh16) : $signed(_GEN_27209); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27211 = 12'h65f == _T_837 ? $signed(7'sh17) : $signed(_GEN_27210); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27212 = 12'h660 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27211); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27213 = 12'h661 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27212); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27214 = 12'h662 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27213); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27215 = 12'h663 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27214); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27216 = 12'h664 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27215); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27217 = 12'h665 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27216); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27218 = 12'h666 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27217); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27219 = 12'h667 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27218); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27220 = 12'h668 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27219); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27221 = 12'h669 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27220); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27222 = 12'h66a == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27221); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27223 = 12'h66b == _T_837 ? $signed(7'sh20) : $signed(_GEN_27222); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27224 = 12'h66c == _T_837 ? $signed(7'sh20) : $signed(_GEN_27223); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27225 = 12'h66d == _T_837 ? $signed(7'sh21) : $signed(_GEN_27224); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27226 = 12'h66e == _T_837 ? $signed(7'sh22) : $signed(_GEN_27225); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27227 = 12'h66f == _T_837 ? $signed(7'sh22) : $signed(_GEN_27226); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27228 = 12'h670 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27227); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27229 = 12'h671 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27228); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27230 = 12'h672 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27229); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27231 = 12'h673 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27230); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27232 = 12'h674 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27231); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27233 = 12'h675 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27232); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27234 = 12'h676 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27233); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27235 = 12'h677 == _T_837 ? $signed(7'sh28) : $signed(_GEN_27234); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27236 = 12'h678 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27235); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27237 = 12'h679 == _T_837 ? $signed(7'sha) : $signed(_GEN_27236); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27238 = 12'h67a == _T_837 ? $signed(7'sha) : $signed(_GEN_27237); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27239 = 12'h67b == _T_837 ? $signed(7'shb) : $signed(_GEN_27238); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27240 = 12'h67c == _T_837 ? $signed(7'shc) : $signed(_GEN_27239); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27241 = 12'h67d == _T_837 ? $signed(7'shc) : $signed(_GEN_27240); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27242 = 12'h67e == _T_837 ? $signed(7'shd) : $signed(_GEN_27241); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27243 = 12'h67f == _T_837 ? $signed(7'she) : $signed(_GEN_27242); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27244 = 12'h680 == _T_837 ? $signed(7'shf) : $signed(_GEN_27243); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27245 = 12'h681 == _T_837 ? $signed(7'shf) : $signed(_GEN_27244); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27246 = 12'h682 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27245); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27247 = 12'h683 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27246); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27248 = 12'h684 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27247); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27249 = 12'h685 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27248); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27250 = 12'h686 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27249); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27251 = 12'h687 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27250); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27252 = 12'h688 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27251); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27253 = 12'h689 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27252); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27254 = 12'h68a == _T_837 ? $signed(7'sh16) : $signed(_GEN_27253); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27255 = 12'h68b == _T_837 ? $signed(7'sh16) : $signed(_GEN_27254); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27256 = 12'h68c == _T_837 ? $signed(7'sh17) : $signed(_GEN_27255); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27257 = 12'h68d == _T_837 ? $signed(7'sh18) : $signed(_GEN_27256); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27258 = 12'h68e == _T_837 ? $signed(7'sh18) : $signed(_GEN_27257); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27259 = 12'h68f == _T_837 ? $signed(7'sh19) : $signed(_GEN_27258); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27260 = 12'h690 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27259); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27261 = 12'h691 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27260); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27262 = 12'h692 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27261); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27263 = 12'h693 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27262); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27264 = 12'h694 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27263); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27265 = 12'h695 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27264); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27266 = 12'h696 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27265); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27267 = 12'h697 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27266); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27268 = 12'h698 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27267); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27269 = 12'h699 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27268); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27270 = 12'h69a == _T_837 ? $signed(7'sh21) : $signed(_GEN_27269); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27271 = 12'h69b == _T_837 ? $signed(7'sh22) : $signed(_GEN_27270); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27272 = 12'h69c == _T_837 ? $signed(7'sh22) : $signed(_GEN_27271); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27273 = 12'h69d == _T_837 ? $signed(7'sh23) : $signed(_GEN_27272); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27274 = 12'h69e == _T_837 ? $signed(7'sh24) : $signed(_GEN_27273); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27275 = 12'h69f == _T_837 ? $signed(7'sh25) : $signed(_GEN_27274); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27276 = 12'h6a0 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27275); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27277 = 12'h6a1 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27276); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27278 = 12'h6a2 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27277); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27279 = 12'h6a3 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27278); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27280 = 12'h6a4 == _T_837 ? $signed(7'sh28) : $signed(_GEN_27279); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27281 = 12'h6a5 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27280); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27282 = 12'h6a6 == _T_837 ? $signed(7'sha) : $signed(_GEN_27281); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27283 = 12'h6a7 == _T_837 ? $signed(7'sha) : $signed(_GEN_27282); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27284 = 12'h6a8 == _T_837 ? $signed(7'shb) : $signed(_GEN_27283); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27285 = 12'h6a9 == _T_837 ? $signed(7'shc) : $signed(_GEN_27284); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27286 = 12'h6aa == _T_837 ? $signed(7'shc) : $signed(_GEN_27285); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27287 = 12'h6ab == _T_837 ? $signed(7'shd) : $signed(_GEN_27286); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27288 = 12'h6ac == _T_837 ? $signed(7'she) : $signed(_GEN_27287); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27289 = 12'h6ad == _T_837 ? $signed(7'shf) : $signed(_GEN_27288); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27290 = 12'h6ae == _T_837 ? $signed(7'shf) : $signed(_GEN_27289); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27291 = 12'h6af == _T_837 ? $signed(7'sh10) : $signed(_GEN_27290); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27292 = 12'h6b0 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27291); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27293 = 12'h6b1 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27292); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27294 = 12'h6b2 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27293); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27295 = 12'h6b3 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27294); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27296 = 12'h6b4 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27295); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27297 = 12'h6b5 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27296); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27298 = 12'h6b6 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27297); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27299 = 12'h6b7 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27298); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27300 = 12'h6b8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27299); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27301 = 12'h6b9 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27300); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27302 = 12'h6ba == _T_837 ? $signed(7'sh18) : $signed(_GEN_27301); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27303 = 12'h6bb == _T_837 ? $signed(7'sh18) : $signed(_GEN_27302); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27304 = 12'h6bc == _T_837 ? $signed(7'sh19) : $signed(_GEN_27303); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27305 = 12'h6bd == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27304); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27306 = 12'h6be == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27305); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27307 = 12'h6bf == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27306); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27308 = 12'h6c0 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27307); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27309 = 12'h6c1 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27308); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27310 = 12'h6c2 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27309); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27311 = 12'h6c3 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27310); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27312 = 12'h6c4 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27311); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27313 = 12'h6c5 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27312); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27314 = 12'h6c6 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27313); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27315 = 12'h6c7 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27314); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27316 = 12'h6c8 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27315); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27317 = 12'h6c9 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27316); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27318 = 12'h6ca == _T_837 ? $signed(7'sh23) : $signed(_GEN_27317); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27319 = 12'h6cb == _T_837 ? $signed(7'sh24) : $signed(_GEN_27318); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27320 = 12'h6cc == _T_837 ? $signed(7'sh25) : $signed(_GEN_27319); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27321 = 12'h6cd == _T_837 ? $signed(7'sh25) : $signed(_GEN_27320); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27322 = 12'h6ce == _T_837 ? $signed(7'sh26) : $signed(_GEN_27321); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27323 = 12'h6cf == _T_837 ? $signed(7'sh27) : $signed(_GEN_27322); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27324 = 12'h6d0 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27323); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27325 = 12'h6d1 == _T_837 ? $signed(7'sh28) : $signed(_GEN_27324); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27326 = 12'h6d2 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27325); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27327 = 12'h6d3 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27326); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27328 = 12'h6d4 == _T_837 ? $signed(7'sha) : $signed(_GEN_27327); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27329 = 12'h6d5 == _T_837 ? $signed(7'shb) : $signed(_GEN_27328); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27330 = 12'h6d6 == _T_837 ? $signed(7'shc) : $signed(_GEN_27329); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27331 = 12'h6d7 == _T_837 ? $signed(7'shc) : $signed(_GEN_27330); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27332 = 12'h6d8 == _T_837 ? $signed(7'shd) : $signed(_GEN_27331); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27333 = 12'h6d9 == _T_837 ? $signed(7'she) : $signed(_GEN_27332); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27334 = 12'h6da == _T_837 ? $signed(7'shf) : $signed(_GEN_27333); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27335 = 12'h6db == _T_837 ? $signed(7'shf) : $signed(_GEN_27334); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27336 = 12'h6dc == _T_837 ? $signed(7'sh10) : $signed(_GEN_27335); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27337 = 12'h6dd == _T_837 ? $signed(7'sh11) : $signed(_GEN_27336); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27338 = 12'h6de == _T_837 ? $signed(7'sh11) : $signed(_GEN_27337); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27339 = 12'h6df == _T_837 ? $signed(7'sh12) : $signed(_GEN_27338); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27340 = 12'h6e0 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27339); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27341 = 12'h6e1 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27340); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27342 = 12'h6e2 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27341); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27343 = 12'h6e3 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27342); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27344 = 12'h6e4 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27343); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27345 = 12'h6e5 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27344); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27346 = 12'h6e6 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27345); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27347 = 12'h6e7 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27346); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27348 = 12'h6e8 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27347); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27349 = 12'h6e9 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27348); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27350 = 12'h6ea == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27349); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27351 = 12'h6eb == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27350); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27352 = 12'h6ec == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27351); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27353 = 12'h6ed == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27352); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27354 = 12'h6ee == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27353); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27355 = 12'h6ef == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27354); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27356 = 12'h6f0 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27355); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27357 = 12'h6f1 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27356); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27358 = 12'h6f2 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27357); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27359 = 12'h6f3 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27358); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27360 = 12'h6f4 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27359); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27361 = 12'h6f5 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27360); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27362 = 12'h6f6 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27361); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27363 = 12'h6f7 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27362); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27364 = 12'h6f8 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27363); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27365 = 12'h6f9 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27364); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27366 = 12'h6fa == _T_837 ? $signed(7'sh25) : $signed(_GEN_27365); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27367 = 12'h6fb == _T_837 ? $signed(7'sh26) : $signed(_GEN_27366); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27368 = 12'h6fc == _T_837 ? $signed(7'sh27) : $signed(_GEN_27367); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27369 = 12'h6fd == _T_837 ? $signed(7'sh27) : $signed(_GEN_27368); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27370 = 12'h6fe == _T_837 ? $signed(7'sh28) : $signed(_GEN_27369); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27371 = 12'h6ff == _T_837 ? $signed(7'sh29) : $signed(_GEN_27370); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27372 = 12'h700 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27371); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27373 = 12'h701 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27372); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27374 = 12'h702 == _T_837 ? $signed(7'shb) : $signed(_GEN_27373); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27375 = 12'h703 == _T_837 ? $signed(7'shc) : $signed(_GEN_27374); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27376 = 12'h704 == _T_837 ? $signed(7'shc) : $signed(_GEN_27375); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27377 = 12'h705 == _T_837 ? $signed(7'shd) : $signed(_GEN_27376); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27378 = 12'h706 == _T_837 ? $signed(7'she) : $signed(_GEN_27377); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27379 = 12'h707 == _T_837 ? $signed(7'shf) : $signed(_GEN_27378); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27380 = 12'h708 == _T_837 ? $signed(7'shf) : $signed(_GEN_27379); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27381 = 12'h709 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27380); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27382 = 12'h70a == _T_837 ? $signed(7'sh11) : $signed(_GEN_27381); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27383 = 12'h70b == _T_837 ? $signed(7'sh11) : $signed(_GEN_27382); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27384 = 12'h70c == _T_837 ? $signed(7'sh12) : $signed(_GEN_27383); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27385 = 12'h70d == _T_837 ? $signed(7'sh13) : $signed(_GEN_27384); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27386 = 12'h70e == _T_837 ? $signed(7'sh14) : $signed(_GEN_27385); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27387 = 12'h70f == _T_837 ? $signed(7'sh14) : $signed(_GEN_27386); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27388 = 12'h710 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27387); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27389 = 12'h711 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27388); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27390 = 12'h712 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27389); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27391 = 12'h713 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27390); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27392 = 12'h714 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27391); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27393 = 12'h715 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27392); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27394 = 12'h716 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27393); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27395 = 12'h717 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27394); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27396 = 12'h718 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27395); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27397 = 12'h719 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27396); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27398 = 12'h71a == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27397); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27399 = 12'h71b == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27398); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27400 = 12'h71c == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27399); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27401 = 12'h71d == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27400); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27402 = 12'h71e == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27401); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27403 = 12'h71f == _T_837 ? $signed(7'sh20) : $signed(_GEN_27402); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27404 = 12'h720 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27403); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27405 = 12'h721 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27404); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27406 = 12'h722 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27405); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27407 = 12'h723 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27406); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27408 = 12'h724 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27407); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27409 = 12'h725 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27408); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27410 = 12'h726 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27409); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27411 = 12'h727 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27410); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27412 = 12'h728 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27411); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27413 = 12'h729 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27412); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27414 = 12'h72a == _T_837 ? $signed(7'sh27) : $signed(_GEN_27413); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27415 = 12'h72b == _T_837 ? $signed(7'sh28) : $signed(_GEN_27414); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27416 = 12'h72c == _T_837 ? $signed(7'sh29) : $signed(_GEN_27415); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27417 = 12'h72d == _T_837 ? $signed(7'sh29) : $signed(_GEN_27416); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27418 = 12'h72e == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27417); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27419 = 12'h72f == _T_837 ? $signed(7'sh2b) : $signed(_GEN_27418); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27420 = 12'h730 == _T_837 ? $signed(7'shc) : $signed(_GEN_27419); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27421 = 12'h731 == _T_837 ? $signed(7'shc) : $signed(_GEN_27420); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27422 = 12'h732 == _T_837 ? $signed(7'shd) : $signed(_GEN_27421); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27423 = 12'h733 == _T_837 ? $signed(7'she) : $signed(_GEN_27422); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27424 = 12'h734 == _T_837 ? $signed(7'shf) : $signed(_GEN_27423); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27425 = 12'h735 == _T_837 ? $signed(7'shf) : $signed(_GEN_27424); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27426 = 12'h736 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27425); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27427 = 12'h737 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27426); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27428 = 12'h738 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27427); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27429 = 12'h739 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27428); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27430 = 12'h73a == _T_837 ? $signed(7'sh13) : $signed(_GEN_27429); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27431 = 12'h73b == _T_837 ? $signed(7'sh14) : $signed(_GEN_27430); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27432 = 12'h73c == _T_837 ? $signed(7'sh14) : $signed(_GEN_27431); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27433 = 12'h73d == _T_837 ? $signed(7'sh15) : $signed(_GEN_27432); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27434 = 12'h73e == _T_837 ? $signed(7'sh16) : $signed(_GEN_27433); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27435 = 12'h73f == _T_837 ? $signed(7'sh16) : $signed(_GEN_27434); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27436 = 12'h740 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27435); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27437 = 12'h741 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27436); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27438 = 12'h742 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27437); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27439 = 12'h743 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27438); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27440 = 12'h744 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27439); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27441 = 12'h745 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27440); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27442 = 12'h746 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27441); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27443 = 12'h747 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27442); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27444 = 12'h748 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27443); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27445 = 12'h749 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27444); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27446 = 12'h74a == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27445); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27447 = 12'h74b == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27446); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27448 = 12'h74c == _T_837 ? $signed(7'sh20) : $signed(_GEN_27447); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27449 = 12'h74d == _T_837 ? $signed(7'sh20) : $signed(_GEN_27448); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27450 = 12'h74e == _T_837 ? $signed(7'sh21) : $signed(_GEN_27449); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27451 = 12'h74f == _T_837 ? $signed(7'sh22) : $signed(_GEN_27450); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27452 = 12'h750 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27451); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27453 = 12'h751 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27452); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27454 = 12'h752 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27453); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27455 = 12'h753 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27454); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27456 = 12'h754 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27455); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27457 = 12'h755 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27456); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27458 = 12'h756 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27457); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27459 = 12'h757 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27458); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27460 = 12'h758 == _T_837 ? $signed(7'sh28) : $signed(_GEN_27459); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27461 = 12'h759 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27460); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27462 = 12'h75a == _T_837 ? $signed(7'sh29) : $signed(_GEN_27461); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27463 = 12'h75b == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27462); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27464 = 12'h75c == _T_837 ? $signed(7'sh2b) : $signed(_GEN_27463); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27465 = 12'h75d == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27464); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27466 = 12'h75e == _T_837 ? $signed(7'shc) : $signed(_GEN_27465); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27467 = 12'h75f == _T_837 ? $signed(7'shd) : $signed(_GEN_27466); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27468 = 12'h760 == _T_837 ? $signed(7'she) : $signed(_GEN_27467); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27469 = 12'h761 == _T_837 ? $signed(7'shf) : $signed(_GEN_27468); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27470 = 12'h762 == _T_837 ? $signed(7'shf) : $signed(_GEN_27469); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27471 = 12'h763 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27470); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27472 = 12'h764 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27471); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27473 = 12'h765 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27472); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27474 = 12'h766 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27473); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27475 = 12'h767 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27474); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27476 = 12'h768 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27475); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27477 = 12'h769 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27476); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27478 = 12'h76a == _T_837 ? $signed(7'sh15) : $signed(_GEN_27477); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27479 = 12'h76b == _T_837 ? $signed(7'sh16) : $signed(_GEN_27478); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27480 = 12'h76c == _T_837 ? $signed(7'sh16) : $signed(_GEN_27479); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27481 = 12'h76d == _T_837 ? $signed(7'sh17) : $signed(_GEN_27480); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27482 = 12'h76e == _T_837 ? $signed(7'sh18) : $signed(_GEN_27481); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27483 = 12'h76f == _T_837 ? $signed(7'sh18) : $signed(_GEN_27482); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27484 = 12'h770 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27483); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27485 = 12'h771 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27484); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27486 = 12'h772 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27485); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27487 = 12'h773 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27486); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27488 = 12'h774 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27487); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27489 = 12'h775 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27488); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27490 = 12'h776 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27489); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27491 = 12'h777 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27490); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27492 = 12'h778 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27491); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27493 = 12'h779 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27492); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27494 = 12'h77a == _T_837 ? $signed(7'sh20) : $signed(_GEN_27493); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27495 = 12'h77b == _T_837 ? $signed(7'sh21) : $signed(_GEN_27494); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27496 = 12'h77c == _T_837 ? $signed(7'sh22) : $signed(_GEN_27495); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27497 = 12'h77d == _T_837 ? $signed(7'sh22) : $signed(_GEN_27496); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27498 = 12'h77e == _T_837 ? $signed(7'sh23) : $signed(_GEN_27497); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27499 = 12'h77f == _T_837 ? $signed(7'sh24) : $signed(_GEN_27498); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27500 = 12'h780 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27499); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27501 = 12'h781 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27500); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27502 = 12'h782 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27501); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27503 = 12'h783 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27502); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27504 = 12'h784 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27503); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27505 = 12'h785 == _T_837 ? $signed(7'sh28) : $signed(_GEN_27504); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27506 = 12'h786 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27505); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27507 = 12'h787 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27506); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27508 = 12'h788 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27507); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27509 = 12'h789 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_27508); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27510 = 12'h78a == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27509); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27511 = 12'h78b == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27510); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27512 = 12'h78c == _T_837 ? $signed(7'shd) : $signed(_GEN_27511); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27513 = 12'h78d == _T_837 ? $signed(7'she) : $signed(_GEN_27512); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27514 = 12'h78e == _T_837 ? $signed(7'shf) : $signed(_GEN_27513); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27515 = 12'h78f == _T_837 ? $signed(7'shf) : $signed(_GEN_27514); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27516 = 12'h790 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27515); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27517 = 12'h791 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27516); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27518 = 12'h792 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27517); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27519 = 12'h793 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27518); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27520 = 12'h794 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27519); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27521 = 12'h795 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27520); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27522 = 12'h796 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27521); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27523 = 12'h797 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27522); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27524 = 12'h798 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27523); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27525 = 12'h799 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27524); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27526 = 12'h79a == _T_837 ? $signed(7'sh17) : $signed(_GEN_27525); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27527 = 12'h79b == _T_837 ? $signed(7'sh18) : $signed(_GEN_27526); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27528 = 12'h79c == _T_837 ? $signed(7'sh18) : $signed(_GEN_27527); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27529 = 12'h79d == _T_837 ? $signed(7'sh19) : $signed(_GEN_27528); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27530 = 12'h79e == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27529); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27531 = 12'h79f == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27530); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27532 = 12'h7a0 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27531); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27533 = 12'h7a1 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27532); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27534 = 12'h7a2 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27533); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27535 = 12'h7a3 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27534); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27536 = 12'h7a4 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27535); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27537 = 12'h7a5 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27536); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27538 = 12'h7a6 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27537); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27539 = 12'h7a7 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27538); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27540 = 12'h7a8 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27539); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27541 = 12'h7a9 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27540); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27542 = 12'h7aa == _T_837 ? $signed(7'sh22) : $signed(_GEN_27541); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27543 = 12'h7ab == _T_837 ? $signed(7'sh23) : $signed(_GEN_27542); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27544 = 12'h7ac == _T_837 ? $signed(7'sh24) : $signed(_GEN_27543); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27545 = 12'h7ad == _T_837 ? $signed(7'sh25) : $signed(_GEN_27544); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27546 = 12'h7ae == _T_837 ? $signed(7'sh25) : $signed(_GEN_27545); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27547 = 12'h7af == _T_837 ? $signed(7'sh26) : $signed(_GEN_27546); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27548 = 12'h7b0 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27547); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27549 = 12'h7b1 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27548); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27550 = 12'h7b2 == _T_837 ? $signed(7'sh28) : $signed(_GEN_27549); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27551 = 12'h7b3 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27550); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27552 = 12'h7b4 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27551); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27553 = 12'h7b5 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27552); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27554 = 12'h7b6 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_27553); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27555 = 12'h7b7 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27554); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27556 = 12'h7b8 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27555); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27557 = 12'h7b9 == _T_837 ? $signed(7'sh2d) : $signed(_GEN_27556); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27558 = 12'h7ba == _T_837 ? $signed(7'she) : $signed(_GEN_27557); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27559 = 12'h7bb == _T_837 ? $signed(7'shf) : $signed(_GEN_27558); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27560 = 12'h7bc == _T_837 ? $signed(7'shf) : $signed(_GEN_27559); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27561 = 12'h7bd == _T_837 ? $signed(7'sh10) : $signed(_GEN_27560); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27562 = 12'h7be == _T_837 ? $signed(7'sh11) : $signed(_GEN_27561); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27563 = 12'h7bf == _T_837 ? $signed(7'sh11) : $signed(_GEN_27562); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27564 = 12'h7c0 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27563); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27565 = 12'h7c1 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27564); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27566 = 12'h7c2 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27565); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27567 = 12'h7c3 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27566); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27568 = 12'h7c4 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27567); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27569 = 12'h7c5 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27568); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27570 = 12'h7c6 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27569); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27571 = 12'h7c7 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27570); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27572 = 12'h7c8 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27571); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27573 = 12'h7c9 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27572); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27574 = 12'h7ca == _T_837 ? $signed(7'sh19) : $signed(_GEN_27573); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27575 = 12'h7cb == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27574); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27576 = 12'h7cc == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27575); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27577 = 12'h7cd == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27576); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27578 = 12'h7ce == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27577); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27579 = 12'h7cf == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27578); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27580 = 12'h7d0 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27579); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27581 = 12'h7d1 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27580); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27582 = 12'h7d2 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27581); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27583 = 12'h7d3 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27582); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27584 = 12'h7d4 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27583); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27585 = 12'h7d5 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27584); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27586 = 12'h7d6 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27585); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27587 = 12'h7d7 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27586); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27588 = 12'h7d8 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27587); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27589 = 12'h7d9 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27588); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27590 = 12'h7da == _T_837 ? $signed(7'sh25) : $signed(_GEN_27589); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27591 = 12'h7db == _T_837 ? $signed(7'sh25) : $signed(_GEN_27590); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27592 = 12'h7dc == _T_837 ? $signed(7'sh26) : $signed(_GEN_27591); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27593 = 12'h7dd == _T_837 ? $signed(7'sh27) : $signed(_GEN_27592); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27594 = 12'h7de == _T_837 ? $signed(7'sh27) : $signed(_GEN_27593); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27595 = 12'h7df == _T_837 ? $signed(7'sh28) : $signed(_GEN_27594); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27596 = 12'h7e0 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27595); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27597 = 12'h7e1 == _T_837 ? $signed(7'sh29) : $signed(_GEN_27596); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27598 = 12'h7e2 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27597); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27599 = 12'h7e3 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_27598); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27600 = 12'h7e4 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27599); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27601 = 12'h7e5 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27600); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27602 = 12'h7e6 == _T_837 ? $signed(7'sh2d) : $signed(_GEN_27601); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27603 = 12'h7e7 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_27602); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27604 = 12'h7e8 == _T_837 ? $signed(7'shf) : $signed(_GEN_27603); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27605 = 12'h7e9 == _T_837 ? $signed(7'shf) : $signed(_GEN_27604); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27606 = 12'h7ea == _T_837 ? $signed(7'sh10) : $signed(_GEN_27605); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27607 = 12'h7eb == _T_837 ? $signed(7'sh11) : $signed(_GEN_27606); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27608 = 12'h7ec == _T_837 ? $signed(7'sh11) : $signed(_GEN_27607); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27609 = 12'h7ed == _T_837 ? $signed(7'sh12) : $signed(_GEN_27608); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27610 = 12'h7ee == _T_837 ? $signed(7'sh13) : $signed(_GEN_27609); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27611 = 12'h7ef == _T_837 ? $signed(7'sh14) : $signed(_GEN_27610); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27612 = 12'h7f0 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27611); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27613 = 12'h7f1 == _T_837 ? $signed(7'sh15) : $signed(_GEN_27612); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27614 = 12'h7f2 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27613); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27615 = 12'h7f3 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27614); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27616 = 12'h7f4 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27615); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27617 = 12'h7f5 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27616); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27618 = 12'h7f6 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27617); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27619 = 12'h7f7 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27618); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27620 = 12'h7f8 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27619); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27621 = 12'h7f9 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27620); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27622 = 12'h7fa == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27621); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27623 = 12'h7fb == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27622); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27624 = 12'h7fc == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27623); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27625 = 12'h7fd == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27624); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27626 = 12'h7fe == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27625); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27627 = 12'h7ff == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27626); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27628 = 12'h800 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27627); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27629 = 12'h801 == _T_837 ? $signed(7'sh20) : $signed(_GEN_27628); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27630 = 12'h802 == _T_837 ? $signed(7'sh21) : $signed(_GEN_27629); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27631 = 12'h803 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27630); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27632 = 12'h804 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27631); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27633 = 12'h805 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27632); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27634 = 12'h806 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27633); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27635 = 12'h807 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27634); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27636 = 12'h808 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27635); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27637 = 12'h809 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27636); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27638 = 12'h80a == _T_837 ? $signed(7'sh27) : $signed(_GEN_27637); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27639 = 12'h80b == _T_837 ? $signed(7'sh27) : $signed(_GEN_27638); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27640 = 12'h80c == _T_837 ? $signed(7'sh28) : $signed(_GEN_27639); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27641 = 12'h80d == _T_837 ? $signed(7'sh29) : $signed(_GEN_27640); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27642 = 12'h80e == _T_837 ? $signed(7'sh29) : $signed(_GEN_27641); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27643 = 12'h80f == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27642); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27644 = 12'h810 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_27643); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27645 = 12'h811 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27644); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27646 = 12'h812 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27645); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27647 = 12'h813 == _T_837 ? $signed(7'sh2d) : $signed(_GEN_27646); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27648 = 12'h814 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_27647); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27649 = 12'h815 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_27648); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27650 = 12'h816 == _T_837 ? $signed(7'shf) : $signed(_GEN_27649); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27651 = 12'h817 == _T_837 ? $signed(7'sh10) : $signed(_GEN_27650); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27652 = 12'h818 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27651); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27653 = 12'h819 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27652); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27654 = 12'h81a == _T_837 ? $signed(7'sh12) : $signed(_GEN_27653); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27655 = 12'h81b == _T_837 ? $signed(7'sh13) : $signed(_GEN_27654); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27656 = 12'h81c == _T_837 ? $signed(7'sh14) : $signed(_GEN_27655); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27657 = 12'h81d == _T_837 ? $signed(7'sh14) : $signed(_GEN_27656); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27658 = 12'h81e == _T_837 ? $signed(7'sh15) : $signed(_GEN_27657); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27659 = 12'h81f == _T_837 ? $signed(7'sh16) : $signed(_GEN_27658); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27660 = 12'h820 == _T_837 ? $signed(7'sh16) : $signed(_GEN_27659); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27661 = 12'h821 == _T_837 ? $signed(7'sh17) : $signed(_GEN_27660); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27662 = 12'h822 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27661); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27663 = 12'h823 == _T_837 ? $signed(7'sh18) : $signed(_GEN_27662); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27664 = 12'h824 == _T_837 ? $signed(7'sh19) : $signed(_GEN_27663); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27665 = 12'h825 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_27664); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27666 = 12'h826 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27665); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27667 = 12'h827 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_27666); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27668 = 12'h828 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_27667); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27669 = 12'h829 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27668); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27670 = 12'h82a == _T_837 ? $signed(7'sh1d) : $signed(_GEN_27669); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27671 = 12'h82b == _T_837 ? $signed(7'sh1e) : $signed(_GEN_27670); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27672 = 12'h82c == _T_837 ? $signed(7'sh1f) : $signed(_GEN_27671); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27673 = 12'h82d == _T_837 ? $signed(7'sh20) : $signed(_GEN_27672); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27674 = 12'h82e == _T_837 ? $signed(7'sh20) : $signed(_GEN_27673); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27675 = 12'h82f == _T_837 ? $signed(7'sh21) : $signed(_GEN_27674); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27676 = 12'h830 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27675); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27677 = 12'h831 == _T_837 ? $signed(7'sh22) : $signed(_GEN_27676); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27678 = 12'h832 == _T_837 ? $signed(7'sh23) : $signed(_GEN_27677); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27679 = 12'h833 == _T_837 ? $signed(7'sh24) : $signed(_GEN_27678); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27680 = 12'h834 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27679); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27681 = 12'h835 == _T_837 ? $signed(7'sh25) : $signed(_GEN_27680); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27682 = 12'h836 == _T_837 ? $signed(7'sh26) : $signed(_GEN_27681); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27683 = 12'h837 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27682); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27684 = 12'h838 == _T_837 ? $signed(7'sh27) : $signed(_GEN_27683); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27685 = 12'h839 == _T_837 ? $signed(7'sh28) : $signed(_GEN_27684); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27686 = 12'h83a == _T_837 ? $signed(7'sh29) : $signed(_GEN_27685); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27687 = 12'h83b == _T_837 ? $signed(7'sh29) : $signed(_GEN_27686); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27688 = 12'h83c == _T_837 ? $signed(7'sh2a) : $signed(_GEN_27687); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27689 = 12'h83d == _T_837 ? $signed(7'sh2b) : $signed(_GEN_27688); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27690 = 12'h83e == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27689); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27691 = 12'h83f == _T_837 ? $signed(7'sh2c) : $signed(_GEN_27690); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27692 = 12'h840 == _T_837 ? $signed(7'sh2d) : $signed(_GEN_27691); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27693 = 12'h841 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_27692); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27694 = 12'h842 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_27693); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27695 = 12'h843 == _T_837 ? $signed(7'sh2f) : $signed(_GEN_27694); // @[GraphicEngineVGA.scala 321:24]
  wire [11:0] inSpriteX_6 = spriteRotationReg_6 ? $signed({{5{_GEN_27695[6]}},_GEN_27695}) : $signed(_T_822); // @[GraphicEngineVGA.scala 321:24]
  wire [6:0] _GEN_27697 = 12'h1 == _T_837 ? $signed(7'shf) : $signed(7'sh10); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27698 = 12'h2 == _T_837 ? $signed(7'shf) : $signed(_GEN_27697); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27699 = 12'h3 == _T_837 ? $signed(7'she) : $signed(_GEN_27698); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27700 = 12'h4 == _T_837 ? $signed(7'shd) : $signed(_GEN_27699); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27701 = 12'h5 == _T_837 ? $signed(7'shc) : $signed(_GEN_27700); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27702 = 12'h6 == _T_837 ? $signed(7'shc) : $signed(_GEN_27701); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27703 = 12'h7 == _T_837 ? $signed(7'shb) : $signed(_GEN_27702); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27704 = 12'h8 == _T_837 ? $signed(7'sha) : $signed(_GEN_27703); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27705 = 12'h9 == _T_837 ? $signed(7'sha) : $signed(_GEN_27704); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27706 = 12'ha == _T_837 ? $signed(7'sh9) : $signed(_GEN_27705); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27707 = 12'hb == _T_837 ? $signed(7'sh8) : $signed(_GEN_27706); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27708 = 12'hc == _T_837 ? $signed(7'sh8) : $signed(_GEN_27707); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27709 = 12'hd == _T_837 ? $signed(7'sh7) : $signed(_GEN_27708); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27710 = 12'he == _T_837 ? $signed(7'sh6) : $signed(_GEN_27709); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27711 = 12'hf == _T_837 ? $signed(7'sh5) : $signed(_GEN_27710); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27712 = 12'h10 == _T_837 ? $signed(7'sh5) : $signed(_GEN_27711); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27713 = 12'h11 == _T_837 ? $signed(7'sh4) : $signed(_GEN_27712); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27714 = 12'h12 == _T_837 ? $signed(7'sh3) : $signed(_GEN_27713); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27715 = 12'h13 == _T_837 ? $signed(7'sh3) : $signed(_GEN_27714); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27716 = 12'h14 == _T_837 ? $signed(7'sh2) : $signed(_GEN_27715); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27717 = 12'h15 == _T_837 ? $signed(7'sh1) : $signed(_GEN_27716); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27718 = 12'h16 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27717); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27719 = 12'h17 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27718); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27720 = 12'h18 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_27719); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27721 = 12'h19 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27720); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27722 = 12'h1a == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27721); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27723 = 12'h1b == _T_837 ? $signed(-7'sh3) : $signed(_GEN_27722); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27724 = 12'h1c == _T_837 ? $signed(-7'sh4) : $signed(_GEN_27723); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27725 = 12'h1d == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27724); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27726 = 12'h1e == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27725); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27727 = 12'h1f == _T_837 ? $signed(-7'sh6) : $signed(_GEN_27726); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27728 = 12'h20 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27727); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27729 = 12'h21 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27728); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27730 = 12'h22 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_27729); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27731 = 12'h23 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27730); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27732 = 12'h24 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27731); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27733 = 12'h25 == _T_837 ? $signed(-7'sha) : $signed(_GEN_27732); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27734 = 12'h26 == _T_837 ? $signed(-7'shb) : $signed(_GEN_27733); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27735 = 12'h27 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27734); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27736 = 12'h28 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27735); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27737 = 12'h29 == _T_837 ? $signed(-7'shd) : $signed(_GEN_27736); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27738 = 12'h2a == _T_837 ? $signed(-7'she) : $signed(_GEN_27737); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27739 = 12'h2b == _T_837 ? $signed(-7'she) : $signed(_GEN_27738); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27740 = 12'h2c == _T_837 ? $signed(-7'shf) : $signed(_GEN_27739); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27741 = 12'h2d == _T_837 ? $signed(-7'sh10) : $signed(_GEN_27740); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27742 = 12'h2e == _T_837 ? $signed(7'sh11) : $signed(_GEN_27741); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27743 = 12'h2f == _T_837 ? $signed(7'sh10) : $signed(_GEN_27742); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27744 = 12'h30 == _T_837 ? $signed(7'shf) : $signed(_GEN_27743); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27745 = 12'h31 == _T_837 ? $signed(7'shf) : $signed(_GEN_27744); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27746 = 12'h32 == _T_837 ? $signed(7'she) : $signed(_GEN_27745); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27747 = 12'h33 == _T_837 ? $signed(7'shd) : $signed(_GEN_27746); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27748 = 12'h34 == _T_837 ? $signed(7'shc) : $signed(_GEN_27747); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27749 = 12'h35 == _T_837 ? $signed(7'shc) : $signed(_GEN_27748); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27750 = 12'h36 == _T_837 ? $signed(7'shb) : $signed(_GEN_27749); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27751 = 12'h37 == _T_837 ? $signed(7'sha) : $signed(_GEN_27750); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27752 = 12'h38 == _T_837 ? $signed(7'sha) : $signed(_GEN_27751); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27753 = 12'h39 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27752); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27754 = 12'h3a == _T_837 ? $signed(7'sh8) : $signed(_GEN_27753); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27755 = 12'h3b == _T_837 ? $signed(7'sh8) : $signed(_GEN_27754); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27756 = 12'h3c == _T_837 ? $signed(7'sh7) : $signed(_GEN_27755); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27757 = 12'h3d == _T_837 ? $signed(7'sh6) : $signed(_GEN_27756); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27758 = 12'h3e == _T_837 ? $signed(7'sh5) : $signed(_GEN_27757); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27759 = 12'h3f == _T_837 ? $signed(7'sh5) : $signed(_GEN_27758); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27760 = 12'h40 == _T_837 ? $signed(7'sh4) : $signed(_GEN_27759); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27761 = 12'h41 == _T_837 ? $signed(7'sh3) : $signed(_GEN_27760); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27762 = 12'h42 == _T_837 ? $signed(7'sh3) : $signed(_GEN_27761); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27763 = 12'h43 == _T_837 ? $signed(7'sh2) : $signed(_GEN_27762); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27764 = 12'h44 == _T_837 ? $signed(7'sh1) : $signed(_GEN_27763); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27765 = 12'h45 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27764); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27766 = 12'h46 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27765); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27767 = 12'h47 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_27766); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27768 = 12'h48 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27767); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27769 = 12'h49 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27768); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27770 = 12'h4a == _T_837 ? $signed(-7'sh3) : $signed(_GEN_27769); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27771 = 12'h4b == _T_837 ? $signed(-7'sh4) : $signed(_GEN_27770); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27772 = 12'h4c == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27771); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27773 = 12'h4d == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27772); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27774 = 12'h4e == _T_837 ? $signed(-7'sh6) : $signed(_GEN_27773); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27775 = 12'h4f == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27774); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27776 = 12'h50 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27775); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27777 = 12'h51 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_27776); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27778 = 12'h52 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27777); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27779 = 12'h53 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27778); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27780 = 12'h54 == _T_837 ? $signed(-7'sha) : $signed(_GEN_27779); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27781 = 12'h55 == _T_837 ? $signed(-7'shb) : $signed(_GEN_27780); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27782 = 12'h56 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27781); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27783 = 12'h57 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27782); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27784 = 12'h58 == _T_837 ? $signed(-7'shd) : $signed(_GEN_27783); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27785 = 12'h59 == _T_837 ? $signed(-7'she) : $signed(_GEN_27784); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27786 = 12'h5a == _T_837 ? $signed(-7'she) : $signed(_GEN_27785); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27787 = 12'h5b == _T_837 ? $signed(-7'shf) : $signed(_GEN_27786); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27788 = 12'h5c == _T_837 ? $signed(7'sh11) : $signed(_GEN_27787); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27789 = 12'h5d == _T_837 ? $signed(7'sh11) : $signed(_GEN_27788); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27790 = 12'h5e == _T_837 ? $signed(7'sh10) : $signed(_GEN_27789); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27791 = 12'h5f == _T_837 ? $signed(7'shf) : $signed(_GEN_27790); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27792 = 12'h60 == _T_837 ? $signed(7'shf) : $signed(_GEN_27791); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27793 = 12'h61 == _T_837 ? $signed(7'she) : $signed(_GEN_27792); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27794 = 12'h62 == _T_837 ? $signed(7'shd) : $signed(_GEN_27793); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27795 = 12'h63 == _T_837 ? $signed(7'shc) : $signed(_GEN_27794); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27796 = 12'h64 == _T_837 ? $signed(7'shc) : $signed(_GEN_27795); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27797 = 12'h65 == _T_837 ? $signed(7'shb) : $signed(_GEN_27796); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27798 = 12'h66 == _T_837 ? $signed(7'sha) : $signed(_GEN_27797); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27799 = 12'h67 == _T_837 ? $signed(7'sha) : $signed(_GEN_27798); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27800 = 12'h68 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27799); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27801 = 12'h69 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27800); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27802 = 12'h6a == _T_837 ? $signed(7'sh8) : $signed(_GEN_27801); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27803 = 12'h6b == _T_837 ? $signed(7'sh7) : $signed(_GEN_27802); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27804 = 12'h6c == _T_837 ? $signed(7'sh6) : $signed(_GEN_27803); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27805 = 12'h6d == _T_837 ? $signed(7'sh5) : $signed(_GEN_27804); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27806 = 12'h6e == _T_837 ? $signed(7'sh5) : $signed(_GEN_27805); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27807 = 12'h6f == _T_837 ? $signed(7'sh4) : $signed(_GEN_27806); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27808 = 12'h70 == _T_837 ? $signed(7'sh3) : $signed(_GEN_27807); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27809 = 12'h71 == _T_837 ? $signed(7'sh3) : $signed(_GEN_27808); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27810 = 12'h72 == _T_837 ? $signed(7'sh2) : $signed(_GEN_27809); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27811 = 12'h73 == _T_837 ? $signed(7'sh1) : $signed(_GEN_27810); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27812 = 12'h74 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27811); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27813 = 12'h75 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27812); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27814 = 12'h76 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_27813); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27815 = 12'h77 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27814); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27816 = 12'h78 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27815); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27817 = 12'h79 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_27816); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27818 = 12'h7a == _T_837 ? $signed(-7'sh4) : $signed(_GEN_27817); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27819 = 12'h7b == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27818); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27820 = 12'h7c == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27819); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27821 = 12'h7d == _T_837 ? $signed(-7'sh6) : $signed(_GEN_27820); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27822 = 12'h7e == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27821); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27823 = 12'h7f == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27822); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27824 = 12'h80 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_27823); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27825 = 12'h81 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27824); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27826 = 12'h82 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27825); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27827 = 12'h83 == _T_837 ? $signed(-7'sha) : $signed(_GEN_27826); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27828 = 12'h84 == _T_837 ? $signed(-7'shb) : $signed(_GEN_27827); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27829 = 12'h85 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27828); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27830 = 12'h86 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27829); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27831 = 12'h87 == _T_837 ? $signed(-7'shd) : $signed(_GEN_27830); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27832 = 12'h88 == _T_837 ? $signed(-7'she) : $signed(_GEN_27831); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27833 = 12'h89 == _T_837 ? $signed(-7'she) : $signed(_GEN_27832); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27834 = 12'h8a == _T_837 ? $signed(7'sh12) : $signed(_GEN_27833); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27835 = 12'h8b == _T_837 ? $signed(7'sh11) : $signed(_GEN_27834); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27836 = 12'h8c == _T_837 ? $signed(7'sh11) : $signed(_GEN_27835); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27837 = 12'h8d == _T_837 ? $signed(7'sh10) : $signed(_GEN_27836); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27838 = 12'h8e == _T_837 ? $signed(7'shf) : $signed(_GEN_27837); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27839 = 12'h8f == _T_837 ? $signed(7'shf) : $signed(_GEN_27838); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27840 = 12'h90 == _T_837 ? $signed(7'she) : $signed(_GEN_27839); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27841 = 12'h91 == _T_837 ? $signed(7'shd) : $signed(_GEN_27840); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27842 = 12'h92 == _T_837 ? $signed(7'shc) : $signed(_GEN_27841); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27843 = 12'h93 == _T_837 ? $signed(7'shc) : $signed(_GEN_27842); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27844 = 12'h94 == _T_837 ? $signed(7'shb) : $signed(_GEN_27843); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27845 = 12'h95 == _T_837 ? $signed(7'sha) : $signed(_GEN_27844); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27846 = 12'h96 == _T_837 ? $signed(7'sha) : $signed(_GEN_27845); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27847 = 12'h97 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27846); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27848 = 12'h98 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27847); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27849 = 12'h99 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27848); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27850 = 12'h9a == _T_837 ? $signed(7'sh7) : $signed(_GEN_27849); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27851 = 12'h9b == _T_837 ? $signed(7'sh6) : $signed(_GEN_27850); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27852 = 12'h9c == _T_837 ? $signed(7'sh5) : $signed(_GEN_27851); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27853 = 12'h9d == _T_837 ? $signed(7'sh5) : $signed(_GEN_27852); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27854 = 12'h9e == _T_837 ? $signed(7'sh4) : $signed(_GEN_27853); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27855 = 12'h9f == _T_837 ? $signed(7'sh3) : $signed(_GEN_27854); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27856 = 12'ha0 == _T_837 ? $signed(7'sh3) : $signed(_GEN_27855); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27857 = 12'ha1 == _T_837 ? $signed(7'sh2) : $signed(_GEN_27856); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27858 = 12'ha2 == _T_837 ? $signed(7'sh1) : $signed(_GEN_27857); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27859 = 12'ha3 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27858); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27860 = 12'ha4 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27859); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27861 = 12'ha5 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_27860); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27862 = 12'ha6 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27861); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27863 = 12'ha7 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27862); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27864 = 12'ha8 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_27863); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27865 = 12'ha9 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_27864); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27866 = 12'haa == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27865); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27867 = 12'hab == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27866); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27868 = 12'hac == _T_837 ? $signed(-7'sh6) : $signed(_GEN_27867); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27869 = 12'had == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27868); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27870 = 12'hae == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27869); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27871 = 12'haf == _T_837 ? $signed(-7'sh8) : $signed(_GEN_27870); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27872 = 12'hb0 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27871); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27873 = 12'hb1 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27872); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27874 = 12'hb2 == _T_837 ? $signed(-7'sha) : $signed(_GEN_27873); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27875 = 12'hb3 == _T_837 ? $signed(-7'shb) : $signed(_GEN_27874); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27876 = 12'hb4 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27875); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27877 = 12'hb5 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27876); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27878 = 12'hb6 == _T_837 ? $signed(-7'shd) : $signed(_GEN_27877); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27879 = 12'hb7 == _T_837 ? $signed(-7'she) : $signed(_GEN_27878); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27880 = 12'hb8 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27879); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27881 = 12'hb9 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27880); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27882 = 12'hba == _T_837 ? $signed(7'sh11) : $signed(_GEN_27881); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27883 = 12'hbb == _T_837 ? $signed(7'sh11) : $signed(_GEN_27882); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27884 = 12'hbc == _T_837 ? $signed(7'sh10) : $signed(_GEN_27883); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27885 = 12'hbd == _T_837 ? $signed(7'shf) : $signed(_GEN_27884); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27886 = 12'hbe == _T_837 ? $signed(7'shf) : $signed(_GEN_27885); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27887 = 12'hbf == _T_837 ? $signed(7'she) : $signed(_GEN_27886); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27888 = 12'hc0 == _T_837 ? $signed(7'shd) : $signed(_GEN_27887); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27889 = 12'hc1 == _T_837 ? $signed(7'shc) : $signed(_GEN_27888); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27890 = 12'hc2 == _T_837 ? $signed(7'shc) : $signed(_GEN_27889); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27891 = 12'hc3 == _T_837 ? $signed(7'shb) : $signed(_GEN_27890); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27892 = 12'hc4 == _T_837 ? $signed(7'sha) : $signed(_GEN_27891); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27893 = 12'hc5 == _T_837 ? $signed(7'sha) : $signed(_GEN_27892); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27894 = 12'hc6 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27893); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27895 = 12'hc7 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27894); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27896 = 12'hc8 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27895); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27897 = 12'hc9 == _T_837 ? $signed(7'sh7) : $signed(_GEN_27896); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27898 = 12'hca == _T_837 ? $signed(7'sh6) : $signed(_GEN_27897); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27899 = 12'hcb == _T_837 ? $signed(7'sh5) : $signed(_GEN_27898); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27900 = 12'hcc == _T_837 ? $signed(7'sh5) : $signed(_GEN_27899); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27901 = 12'hcd == _T_837 ? $signed(7'sh4) : $signed(_GEN_27900); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27902 = 12'hce == _T_837 ? $signed(7'sh3) : $signed(_GEN_27901); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27903 = 12'hcf == _T_837 ? $signed(7'sh3) : $signed(_GEN_27902); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27904 = 12'hd0 == _T_837 ? $signed(7'sh2) : $signed(_GEN_27903); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27905 = 12'hd1 == _T_837 ? $signed(7'sh1) : $signed(_GEN_27904); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27906 = 12'hd2 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27905); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27907 = 12'hd3 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27906); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27908 = 12'hd4 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_27907); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27909 = 12'hd5 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27908); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27910 = 12'hd6 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27909); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27911 = 12'hd7 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_27910); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27912 = 12'hd8 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_27911); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27913 = 12'hd9 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27912); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27914 = 12'hda == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27913); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27915 = 12'hdb == _T_837 ? $signed(-7'sh6) : $signed(_GEN_27914); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27916 = 12'hdc == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27915); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27917 = 12'hdd == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27916); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27918 = 12'hde == _T_837 ? $signed(-7'sh8) : $signed(_GEN_27917); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27919 = 12'hdf == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27918); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27920 = 12'he0 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27919); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27921 = 12'he1 == _T_837 ? $signed(-7'sha) : $signed(_GEN_27920); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27922 = 12'he2 == _T_837 ? $signed(-7'shb) : $signed(_GEN_27921); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27923 = 12'he3 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27922); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27924 = 12'he4 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27923); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27925 = 12'he5 == _T_837 ? $signed(-7'shd) : $signed(_GEN_27924); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27926 = 12'he6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27925); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27927 = 12'he7 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27926); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27928 = 12'he8 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27927); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27929 = 12'he9 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27928); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27930 = 12'hea == _T_837 ? $signed(7'sh11) : $signed(_GEN_27929); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27931 = 12'heb == _T_837 ? $signed(7'sh10) : $signed(_GEN_27930); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27932 = 12'hec == _T_837 ? $signed(7'shf) : $signed(_GEN_27931); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27933 = 12'hed == _T_837 ? $signed(7'shf) : $signed(_GEN_27932); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27934 = 12'hee == _T_837 ? $signed(7'she) : $signed(_GEN_27933); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27935 = 12'hef == _T_837 ? $signed(7'shd) : $signed(_GEN_27934); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27936 = 12'hf0 == _T_837 ? $signed(7'shc) : $signed(_GEN_27935); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27937 = 12'hf1 == _T_837 ? $signed(7'shc) : $signed(_GEN_27936); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27938 = 12'hf2 == _T_837 ? $signed(7'shb) : $signed(_GEN_27937); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27939 = 12'hf3 == _T_837 ? $signed(7'sha) : $signed(_GEN_27938); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27940 = 12'hf4 == _T_837 ? $signed(7'sha) : $signed(_GEN_27939); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27941 = 12'hf5 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27940); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27942 = 12'hf6 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27941); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27943 = 12'hf7 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27942); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27944 = 12'hf8 == _T_837 ? $signed(7'sh7) : $signed(_GEN_27943); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27945 = 12'hf9 == _T_837 ? $signed(7'sh6) : $signed(_GEN_27944); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27946 = 12'hfa == _T_837 ? $signed(7'sh5) : $signed(_GEN_27945); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27947 = 12'hfb == _T_837 ? $signed(7'sh5) : $signed(_GEN_27946); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27948 = 12'hfc == _T_837 ? $signed(7'sh4) : $signed(_GEN_27947); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27949 = 12'hfd == _T_837 ? $signed(7'sh3) : $signed(_GEN_27948); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27950 = 12'hfe == _T_837 ? $signed(7'sh3) : $signed(_GEN_27949); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27951 = 12'hff == _T_837 ? $signed(7'sh2) : $signed(_GEN_27950); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27952 = 12'h100 == _T_837 ? $signed(7'sh1) : $signed(_GEN_27951); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27953 = 12'h101 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27952); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27954 = 12'h102 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27953); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27955 = 12'h103 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_27954); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27956 = 12'h104 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27955); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27957 = 12'h105 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_27956); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27958 = 12'h106 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_27957); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27959 = 12'h107 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_27958); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27960 = 12'h108 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27959); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27961 = 12'h109 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_27960); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27962 = 12'h10a == _T_837 ? $signed(-7'sh6) : $signed(_GEN_27961); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27963 = 12'h10b == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27962); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27964 = 12'h10c == _T_837 ? $signed(-7'sh7) : $signed(_GEN_27963); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27965 = 12'h10d == _T_837 ? $signed(-7'sh8) : $signed(_GEN_27964); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27966 = 12'h10e == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27965); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27967 = 12'h10f == _T_837 ? $signed(-7'sh9) : $signed(_GEN_27966); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27968 = 12'h110 == _T_837 ? $signed(-7'sha) : $signed(_GEN_27967); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27969 = 12'h111 == _T_837 ? $signed(-7'shb) : $signed(_GEN_27968); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27970 = 12'h112 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27969); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27971 = 12'h113 == _T_837 ? $signed(-7'shc) : $signed(_GEN_27970); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27972 = 12'h114 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27971); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27973 = 12'h115 == _T_837 ? $signed(7'sh14) : $signed(_GEN_27972); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27974 = 12'h116 == _T_837 ? $signed(7'sh13) : $signed(_GEN_27973); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27975 = 12'h117 == _T_837 ? $signed(7'sh12) : $signed(_GEN_27974); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27976 = 12'h118 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27975); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27977 = 12'h119 == _T_837 ? $signed(7'sh11) : $signed(_GEN_27976); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27978 = 12'h11a == _T_837 ? $signed(7'sh10) : $signed(_GEN_27977); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27979 = 12'h11b == _T_837 ? $signed(7'shf) : $signed(_GEN_27978); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27980 = 12'h11c == _T_837 ? $signed(7'shf) : $signed(_GEN_27979); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27981 = 12'h11d == _T_837 ? $signed(7'she) : $signed(_GEN_27980); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27982 = 12'h11e == _T_837 ? $signed(7'shd) : $signed(_GEN_27981); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27983 = 12'h11f == _T_837 ? $signed(7'shc) : $signed(_GEN_27982); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27984 = 12'h120 == _T_837 ? $signed(7'shc) : $signed(_GEN_27983); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27985 = 12'h121 == _T_837 ? $signed(7'shb) : $signed(_GEN_27984); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27986 = 12'h122 == _T_837 ? $signed(7'sha) : $signed(_GEN_27985); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27987 = 12'h123 == _T_837 ? $signed(7'sha) : $signed(_GEN_27986); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27988 = 12'h124 == _T_837 ? $signed(7'sh9) : $signed(_GEN_27987); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27989 = 12'h125 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27988); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27990 = 12'h126 == _T_837 ? $signed(7'sh8) : $signed(_GEN_27989); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27991 = 12'h127 == _T_837 ? $signed(7'sh7) : $signed(_GEN_27990); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27992 = 12'h128 == _T_837 ? $signed(7'sh6) : $signed(_GEN_27991); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27993 = 12'h129 == _T_837 ? $signed(7'sh5) : $signed(_GEN_27992); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27994 = 12'h12a == _T_837 ? $signed(7'sh5) : $signed(_GEN_27993); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27995 = 12'h12b == _T_837 ? $signed(7'sh4) : $signed(_GEN_27994); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27996 = 12'h12c == _T_837 ? $signed(7'sh3) : $signed(_GEN_27995); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27997 = 12'h12d == _T_837 ? $signed(7'sh3) : $signed(_GEN_27996); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27998 = 12'h12e == _T_837 ? $signed(7'sh2) : $signed(_GEN_27997); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_27999 = 12'h12f == _T_837 ? $signed(7'sh1) : $signed(_GEN_27998); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28000 = 12'h130 == _T_837 ? $signed(7'sh0) : $signed(_GEN_27999); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28001 = 12'h131 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28000); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28002 = 12'h132 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28001); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28003 = 12'h133 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28002); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28004 = 12'h134 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28003); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28005 = 12'h135 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28004); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28006 = 12'h136 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28005); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28007 = 12'h137 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28006); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28008 = 12'h138 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28007); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28009 = 12'h139 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28008); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28010 = 12'h13a == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28009); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28011 = 12'h13b == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28010); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28012 = 12'h13c == _T_837 ? $signed(-7'sh8) : $signed(_GEN_28011); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28013 = 12'h13d == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28012); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28014 = 12'h13e == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28013); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28015 = 12'h13f == _T_837 ? $signed(-7'sha) : $signed(_GEN_28014); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28016 = 12'h140 == _T_837 ? $signed(-7'shb) : $signed(_GEN_28015); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28017 = 12'h141 == _T_837 ? $signed(-7'shc) : $signed(_GEN_28016); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28018 = 12'h142 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28017); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28019 = 12'h143 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28018); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28020 = 12'h144 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28019); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28021 = 12'h145 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28020); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28022 = 12'h146 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28021); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28023 = 12'h147 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28022); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28024 = 12'h148 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28023); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28025 = 12'h149 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28024); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28026 = 12'h14a == _T_837 ? $signed(7'shf) : $signed(_GEN_28025); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28027 = 12'h14b == _T_837 ? $signed(7'shf) : $signed(_GEN_28026); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28028 = 12'h14c == _T_837 ? $signed(7'she) : $signed(_GEN_28027); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28029 = 12'h14d == _T_837 ? $signed(7'shd) : $signed(_GEN_28028); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28030 = 12'h14e == _T_837 ? $signed(7'shc) : $signed(_GEN_28029); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28031 = 12'h14f == _T_837 ? $signed(7'shc) : $signed(_GEN_28030); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28032 = 12'h150 == _T_837 ? $signed(7'shb) : $signed(_GEN_28031); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28033 = 12'h151 == _T_837 ? $signed(7'sha) : $signed(_GEN_28032); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28034 = 12'h152 == _T_837 ? $signed(7'sha) : $signed(_GEN_28033); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28035 = 12'h153 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28034); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28036 = 12'h154 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28035); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28037 = 12'h155 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28036); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28038 = 12'h156 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28037); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28039 = 12'h157 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28038); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28040 = 12'h158 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28039); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28041 = 12'h159 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28040); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28042 = 12'h15a == _T_837 ? $signed(7'sh4) : $signed(_GEN_28041); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28043 = 12'h15b == _T_837 ? $signed(7'sh3) : $signed(_GEN_28042); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28044 = 12'h15c == _T_837 ? $signed(7'sh3) : $signed(_GEN_28043); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28045 = 12'h15d == _T_837 ? $signed(7'sh2) : $signed(_GEN_28044); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28046 = 12'h15e == _T_837 ? $signed(7'sh1) : $signed(_GEN_28045); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28047 = 12'h15f == _T_837 ? $signed(7'sh0) : $signed(_GEN_28046); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28048 = 12'h160 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28047); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28049 = 12'h161 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28048); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28050 = 12'h162 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28049); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28051 = 12'h163 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28050); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28052 = 12'h164 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28051); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28053 = 12'h165 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28052); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28054 = 12'h166 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28053); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28055 = 12'h167 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28054); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28056 = 12'h168 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28055); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28057 = 12'h169 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28056); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28058 = 12'h16a == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28057); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28059 = 12'h16b == _T_837 ? $signed(-7'sh8) : $signed(_GEN_28058); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28060 = 12'h16c == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28059); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28061 = 12'h16d == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28060); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28062 = 12'h16e == _T_837 ? $signed(-7'sha) : $signed(_GEN_28061); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28063 = 12'h16f == _T_837 ? $signed(-7'shb) : $signed(_GEN_28062); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28064 = 12'h170 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28063); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28065 = 12'h171 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28064); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28066 = 12'h172 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28065); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28067 = 12'h173 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28066); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28068 = 12'h174 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28067); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28069 = 12'h175 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28068); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28070 = 12'h176 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28069); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28071 = 12'h177 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28070); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28072 = 12'h178 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28071); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28073 = 12'h179 == _T_837 ? $signed(7'shf) : $signed(_GEN_28072); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28074 = 12'h17a == _T_837 ? $signed(7'shf) : $signed(_GEN_28073); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28075 = 12'h17b == _T_837 ? $signed(7'she) : $signed(_GEN_28074); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28076 = 12'h17c == _T_837 ? $signed(7'shd) : $signed(_GEN_28075); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28077 = 12'h17d == _T_837 ? $signed(7'shc) : $signed(_GEN_28076); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28078 = 12'h17e == _T_837 ? $signed(7'shc) : $signed(_GEN_28077); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28079 = 12'h17f == _T_837 ? $signed(7'shb) : $signed(_GEN_28078); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28080 = 12'h180 == _T_837 ? $signed(7'sha) : $signed(_GEN_28079); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28081 = 12'h181 == _T_837 ? $signed(7'sha) : $signed(_GEN_28080); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28082 = 12'h182 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28081); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28083 = 12'h183 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28082); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28084 = 12'h184 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28083); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28085 = 12'h185 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28084); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28086 = 12'h186 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28085); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28087 = 12'h187 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28086); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28088 = 12'h188 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28087); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28089 = 12'h189 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28088); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28090 = 12'h18a == _T_837 ? $signed(7'sh3) : $signed(_GEN_28089); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28091 = 12'h18b == _T_837 ? $signed(7'sh3) : $signed(_GEN_28090); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28092 = 12'h18c == _T_837 ? $signed(7'sh2) : $signed(_GEN_28091); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28093 = 12'h18d == _T_837 ? $signed(7'sh1) : $signed(_GEN_28092); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28094 = 12'h18e == _T_837 ? $signed(7'sh0) : $signed(_GEN_28093); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28095 = 12'h18f == _T_837 ? $signed(7'sh0) : $signed(_GEN_28094); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28096 = 12'h190 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28095); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28097 = 12'h191 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28096); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28098 = 12'h192 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28097); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28099 = 12'h193 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28098); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28100 = 12'h194 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28099); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28101 = 12'h195 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28100); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28102 = 12'h196 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28101); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28103 = 12'h197 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28102); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28104 = 12'h198 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28103); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28105 = 12'h199 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28104); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28106 = 12'h19a == _T_837 ? $signed(-7'sh8) : $signed(_GEN_28105); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28107 = 12'h19b == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28106); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28108 = 12'h19c == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28107); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28109 = 12'h19d == _T_837 ? $signed(-7'sha) : $signed(_GEN_28108); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28110 = 12'h19e == _T_837 ? $signed(7'sh16) : $signed(_GEN_28109); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28111 = 12'h19f == _T_837 ? $signed(7'sh16) : $signed(_GEN_28110); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28112 = 12'h1a0 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28111); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28113 = 12'h1a1 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28112); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28114 = 12'h1a2 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28113); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28115 = 12'h1a3 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28114); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28116 = 12'h1a4 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28115); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28117 = 12'h1a5 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28116); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28118 = 12'h1a6 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28117); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28119 = 12'h1a7 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28118); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28120 = 12'h1a8 == _T_837 ? $signed(7'shf) : $signed(_GEN_28119); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28121 = 12'h1a9 == _T_837 ? $signed(7'shf) : $signed(_GEN_28120); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28122 = 12'h1aa == _T_837 ? $signed(7'she) : $signed(_GEN_28121); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28123 = 12'h1ab == _T_837 ? $signed(7'shd) : $signed(_GEN_28122); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28124 = 12'h1ac == _T_837 ? $signed(7'shc) : $signed(_GEN_28123); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28125 = 12'h1ad == _T_837 ? $signed(7'shc) : $signed(_GEN_28124); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28126 = 12'h1ae == _T_837 ? $signed(7'shb) : $signed(_GEN_28125); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28127 = 12'h1af == _T_837 ? $signed(7'sha) : $signed(_GEN_28126); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28128 = 12'h1b0 == _T_837 ? $signed(7'sha) : $signed(_GEN_28127); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28129 = 12'h1b1 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28128); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28130 = 12'h1b2 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28129); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28131 = 12'h1b3 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28130); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28132 = 12'h1b4 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28131); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28133 = 12'h1b5 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28132); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28134 = 12'h1b6 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28133); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28135 = 12'h1b7 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28134); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28136 = 12'h1b8 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28135); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28137 = 12'h1b9 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28136); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28138 = 12'h1ba == _T_837 ? $signed(7'sh3) : $signed(_GEN_28137); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28139 = 12'h1bb == _T_837 ? $signed(7'sh2) : $signed(_GEN_28138); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28140 = 12'h1bc == _T_837 ? $signed(7'sh1) : $signed(_GEN_28139); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28141 = 12'h1bd == _T_837 ? $signed(7'sh0) : $signed(_GEN_28140); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28142 = 12'h1be == _T_837 ? $signed(7'sh0) : $signed(_GEN_28141); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28143 = 12'h1bf == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28142); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28144 = 12'h1c0 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28143); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28145 = 12'h1c1 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28144); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28146 = 12'h1c2 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28145); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28147 = 12'h1c3 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28146); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28148 = 12'h1c4 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28147); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28149 = 12'h1c5 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28148); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28150 = 12'h1c6 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28149); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28151 = 12'h1c7 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28150); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28152 = 12'h1c8 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28151); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28153 = 12'h1c9 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_28152); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28154 = 12'h1ca == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28153); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28155 = 12'h1cb == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28154); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28156 = 12'h1cc == _T_837 ? $signed(7'sh17) : $signed(_GEN_28155); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28157 = 12'h1cd == _T_837 ? $signed(7'sh16) : $signed(_GEN_28156); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28158 = 12'h1ce == _T_837 ? $signed(7'sh16) : $signed(_GEN_28157); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28159 = 12'h1cf == _T_837 ? $signed(7'sh15) : $signed(_GEN_28158); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28160 = 12'h1d0 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28159); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28161 = 12'h1d1 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28160); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28162 = 12'h1d2 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28161); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28163 = 12'h1d3 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28162); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28164 = 12'h1d4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28163); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28165 = 12'h1d5 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28164); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28166 = 12'h1d6 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28165); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28167 = 12'h1d7 == _T_837 ? $signed(7'shf) : $signed(_GEN_28166); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28168 = 12'h1d8 == _T_837 ? $signed(7'shf) : $signed(_GEN_28167); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28169 = 12'h1d9 == _T_837 ? $signed(7'she) : $signed(_GEN_28168); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28170 = 12'h1da == _T_837 ? $signed(7'shd) : $signed(_GEN_28169); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28171 = 12'h1db == _T_837 ? $signed(7'shc) : $signed(_GEN_28170); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28172 = 12'h1dc == _T_837 ? $signed(7'shc) : $signed(_GEN_28171); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28173 = 12'h1dd == _T_837 ? $signed(7'shb) : $signed(_GEN_28172); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28174 = 12'h1de == _T_837 ? $signed(7'sha) : $signed(_GEN_28173); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28175 = 12'h1df == _T_837 ? $signed(7'sha) : $signed(_GEN_28174); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28176 = 12'h1e0 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28175); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28177 = 12'h1e1 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28176); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28178 = 12'h1e2 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28177); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28179 = 12'h1e3 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28178); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28180 = 12'h1e4 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28179); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28181 = 12'h1e5 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28180); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28182 = 12'h1e6 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28181); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28183 = 12'h1e7 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28182); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28184 = 12'h1e8 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28183); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28185 = 12'h1e9 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28184); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28186 = 12'h1ea == _T_837 ? $signed(7'sh2) : $signed(_GEN_28185); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28187 = 12'h1eb == _T_837 ? $signed(7'sh1) : $signed(_GEN_28186); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28188 = 12'h1ec == _T_837 ? $signed(7'sh0) : $signed(_GEN_28187); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28189 = 12'h1ed == _T_837 ? $signed(7'sh0) : $signed(_GEN_28188); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28190 = 12'h1ee == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28189); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28191 = 12'h1ef == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28190); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28192 = 12'h1f0 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28191); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28193 = 12'h1f1 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28192); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28194 = 12'h1f2 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28193); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28195 = 12'h1f3 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28194); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28196 = 12'h1f4 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28195); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28197 = 12'h1f5 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28196); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28198 = 12'h1f6 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28197); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28199 = 12'h1f7 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28198); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28200 = 12'h1f8 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_28199); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28201 = 12'h1f9 == _T_837 ? $signed(-7'sh9) : $signed(_GEN_28200); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28202 = 12'h1fa == _T_837 ? $signed(7'sh18) : $signed(_GEN_28201); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28203 = 12'h1fb == _T_837 ? $signed(7'sh17) : $signed(_GEN_28202); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28204 = 12'h1fc == _T_837 ? $signed(7'sh16) : $signed(_GEN_28203); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28205 = 12'h1fd == _T_837 ? $signed(7'sh16) : $signed(_GEN_28204); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28206 = 12'h1fe == _T_837 ? $signed(7'sh15) : $signed(_GEN_28205); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28207 = 12'h1ff == _T_837 ? $signed(7'sh14) : $signed(_GEN_28206); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28208 = 12'h200 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28207); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28209 = 12'h201 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28208); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28210 = 12'h202 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28209); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28211 = 12'h203 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28210); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28212 = 12'h204 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28211); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28213 = 12'h205 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28212); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28214 = 12'h206 == _T_837 ? $signed(7'shf) : $signed(_GEN_28213); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28215 = 12'h207 == _T_837 ? $signed(7'shf) : $signed(_GEN_28214); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28216 = 12'h208 == _T_837 ? $signed(7'she) : $signed(_GEN_28215); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28217 = 12'h209 == _T_837 ? $signed(7'shd) : $signed(_GEN_28216); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28218 = 12'h20a == _T_837 ? $signed(7'shc) : $signed(_GEN_28217); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28219 = 12'h20b == _T_837 ? $signed(7'shc) : $signed(_GEN_28218); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28220 = 12'h20c == _T_837 ? $signed(7'shb) : $signed(_GEN_28219); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28221 = 12'h20d == _T_837 ? $signed(7'sha) : $signed(_GEN_28220); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28222 = 12'h20e == _T_837 ? $signed(7'sha) : $signed(_GEN_28221); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28223 = 12'h20f == _T_837 ? $signed(7'sh9) : $signed(_GEN_28222); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28224 = 12'h210 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28223); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28225 = 12'h211 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28224); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28226 = 12'h212 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28225); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28227 = 12'h213 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28226); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28228 = 12'h214 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28227); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28229 = 12'h215 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28228); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28230 = 12'h216 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28229); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28231 = 12'h217 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28230); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28232 = 12'h218 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28231); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28233 = 12'h219 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28232); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28234 = 12'h21a == _T_837 ? $signed(7'sh1) : $signed(_GEN_28233); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28235 = 12'h21b == _T_837 ? $signed(7'sh0) : $signed(_GEN_28234); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28236 = 12'h21c == _T_837 ? $signed(7'sh0) : $signed(_GEN_28235); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28237 = 12'h21d == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28236); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28238 = 12'h21e == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28237); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28239 = 12'h21f == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28238); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28240 = 12'h220 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28239); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28241 = 12'h221 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28240); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28242 = 12'h222 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28241); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28243 = 12'h223 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28242); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28244 = 12'h224 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28243); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28245 = 12'h225 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28244); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28246 = 12'h226 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28245); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28247 = 12'h227 == _T_837 ? $signed(-7'sh8) : $signed(_GEN_28246); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28248 = 12'h228 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28247); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28249 = 12'h229 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28248); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28250 = 12'h22a == _T_837 ? $signed(7'sh17) : $signed(_GEN_28249); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28251 = 12'h22b == _T_837 ? $signed(7'sh16) : $signed(_GEN_28250); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28252 = 12'h22c == _T_837 ? $signed(7'sh16) : $signed(_GEN_28251); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28253 = 12'h22d == _T_837 ? $signed(7'sh15) : $signed(_GEN_28252); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28254 = 12'h22e == _T_837 ? $signed(7'sh14) : $signed(_GEN_28253); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28255 = 12'h22f == _T_837 ? $signed(7'sh14) : $signed(_GEN_28254); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28256 = 12'h230 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28255); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28257 = 12'h231 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28256); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28258 = 12'h232 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28257); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28259 = 12'h233 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28258); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28260 = 12'h234 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28259); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28261 = 12'h235 == _T_837 ? $signed(7'shf) : $signed(_GEN_28260); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28262 = 12'h236 == _T_837 ? $signed(7'shf) : $signed(_GEN_28261); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28263 = 12'h237 == _T_837 ? $signed(7'she) : $signed(_GEN_28262); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28264 = 12'h238 == _T_837 ? $signed(7'shd) : $signed(_GEN_28263); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28265 = 12'h239 == _T_837 ? $signed(7'shc) : $signed(_GEN_28264); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28266 = 12'h23a == _T_837 ? $signed(7'shc) : $signed(_GEN_28265); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28267 = 12'h23b == _T_837 ? $signed(7'shb) : $signed(_GEN_28266); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28268 = 12'h23c == _T_837 ? $signed(7'sha) : $signed(_GEN_28267); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28269 = 12'h23d == _T_837 ? $signed(7'sha) : $signed(_GEN_28268); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28270 = 12'h23e == _T_837 ? $signed(7'sh9) : $signed(_GEN_28269); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28271 = 12'h23f == _T_837 ? $signed(7'sh8) : $signed(_GEN_28270); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28272 = 12'h240 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28271); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28273 = 12'h241 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28272); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28274 = 12'h242 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28273); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28275 = 12'h243 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28274); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28276 = 12'h244 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28275); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28277 = 12'h245 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28276); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28278 = 12'h246 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28277); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28279 = 12'h247 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28278); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28280 = 12'h248 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28279); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28281 = 12'h249 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28280); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28282 = 12'h24a == _T_837 ? $signed(7'sh0) : $signed(_GEN_28281); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28283 = 12'h24b == _T_837 ? $signed(7'sh0) : $signed(_GEN_28282); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28284 = 12'h24c == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28283); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28285 = 12'h24d == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28284); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28286 = 12'h24e == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28285); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28287 = 12'h24f == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28286); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28288 = 12'h250 == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28287); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28289 = 12'h251 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28288); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28290 = 12'h252 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28289); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28291 = 12'h253 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28290); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28292 = 12'h254 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28291); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28293 = 12'h255 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28292); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28294 = 12'h256 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28293); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28295 = 12'h257 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28294); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28296 = 12'h258 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28295); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28297 = 12'h259 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28296); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28298 = 12'h25a == _T_837 ? $signed(7'sh16) : $signed(_GEN_28297); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28299 = 12'h25b == _T_837 ? $signed(7'sh16) : $signed(_GEN_28298); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28300 = 12'h25c == _T_837 ? $signed(7'sh15) : $signed(_GEN_28299); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28301 = 12'h25d == _T_837 ? $signed(7'sh14) : $signed(_GEN_28300); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28302 = 12'h25e == _T_837 ? $signed(7'sh14) : $signed(_GEN_28301); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28303 = 12'h25f == _T_837 ? $signed(7'sh13) : $signed(_GEN_28302); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28304 = 12'h260 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28303); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28305 = 12'h261 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28304); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28306 = 12'h262 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28305); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28307 = 12'h263 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28306); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28308 = 12'h264 == _T_837 ? $signed(7'shf) : $signed(_GEN_28307); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28309 = 12'h265 == _T_837 ? $signed(7'shf) : $signed(_GEN_28308); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28310 = 12'h266 == _T_837 ? $signed(7'she) : $signed(_GEN_28309); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28311 = 12'h267 == _T_837 ? $signed(7'shd) : $signed(_GEN_28310); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28312 = 12'h268 == _T_837 ? $signed(7'shc) : $signed(_GEN_28311); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28313 = 12'h269 == _T_837 ? $signed(7'shc) : $signed(_GEN_28312); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28314 = 12'h26a == _T_837 ? $signed(7'shb) : $signed(_GEN_28313); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28315 = 12'h26b == _T_837 ? $signed(7'sha) : $signed(_GEN_28314); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28316 = 12'h26c == _T_837 ? $signed(7'sha) : $signed(_GEN_28315); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28317 = 12'h26d == _T_837 ? $signed(7'sh9) : $signed(_GEN_28316); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28318 = 12'h26e == _T_837 ? $signed(7'sh8) : $signed(_GEN_28317); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28319 = 12'h26f == _T_837 ? $signed(7'sh8) : $signed(_GEN_28318); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28320 = 12'h270 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28319); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28321 = 12'h271 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28320); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28322 = 12'h272 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28321); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28323 = 12'h273 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28322); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28324 = 12'h274 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28323); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28325 = 12'h275 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28324); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28326 = 12'h276 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28325); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28327 = 12'h277 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28326); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28328 = 12'h278 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28327); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28329 = 12'h279 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28328); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28330 = 12'h27a == _T_837 ? $signed(7'sh0) : $signed(_GEN_28329); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28331 = 12'h27b == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28330); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28332 = 12'h27c == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28331); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28333 = 12'h27d == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28332); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28334 = 12'h27e == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28333); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28335 = 12'h27f == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28334); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28336 = 12'h280 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28335); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28337 = 12'h281 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28336); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28338 = 12'h282 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28337); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28339 = 12'h283 == _T_837 ? $signed(-7'sh7) : $signed(_GEN_28338); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28340 = 12'h284 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28339); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28341 = 12'h285 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28340); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28342 = 12'h286 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28341); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28343 = 12'h287 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28342); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28344 = 12'h288 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28343); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28345 = 12'h289 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28344); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28346 = 12'h28a == _T_837 ? $signed(7'sh16) : $signed(_GEN_28345); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28347 = 12'h28b == _T_837 ? $signed(7'sh15) : $signed(_GEN_28346); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28348 = 12'h28c == _T_837 ? $signed(7'sh14) : $signed(_GEN_28347); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28349 = 12'h28d == _T_837 ? $signed(7'sh14) : $signed(_GEN_28348); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28350 = 12'h28e == _T_837 ? $signed(7'sh13) : $signed(_GEN_28349); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28351 = 12'h28f == _T_837 ? $signed(7'sh12) : $signed(_GEN_28350); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28352 = 12'h290 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28351); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28353 = 12'h291 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28352); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28354 = 12'h292 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28353); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28355 = 12'h293 == _T_837 ? $signed(7'shf) : $signed(_GEN_28354); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28356 = 12'h294 == _T_837 ? $signed(7'shf) : $signed(_GEN_28355); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28357 = 12'h295 == _T_837 ? $signed(7'she) : $signed(_GEN_28356); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28358 = 12'h296 == _T_837 ? $signed(7'shd) : $signed(_GEN_28357); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28359 = 12'h297 == _T_837 ? $signed(7'shc) : $signed(_GEN_28358); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28360 = 12'h298 == _T_837 ? $signed(7'shc) : $signed(_GEN_28359); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28361 = 12'h299 == _T_837 ? $signed(7'shb) : $signed(_GEN_28360); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28362 = 12'h29a == _T_837 ? $signed(7'sha) : $signed(_GEN_28361); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28363 = 12'h29b == _T_837 ? $signed(7'sha) : $signed(_GEN_28362); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28364 = 12'h29c == _T_837 ? $signed(7'sh9) : $signed(_GEN_28363); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28365 = 12'h29d == _T_837 ? $signed(7'sh8) : $signed(_GEN_28364); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28366 = 12'h29e == _T_837 ? $signed(7'sh8) : $signed(_GEN_28365); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28367 = 12'h29f == _T_837 ? $signed(7'sh7) : $signed(_GEN_28366); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28368 = 12'h2a0 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28367); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28369 = 12'h2a1 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28368); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28370 = 12'h2a2 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28369); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28371 = 12'h2a3 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28370); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28372 = 12'h2a4 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28371); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28373 = 12'h2a5 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28372); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28374 = 12'h2a6 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28373); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28375 = 12'h2a7 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28374); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28376 = 12'h2a8 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28375); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28377 = 12'h2a9 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28376); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28378 = 12'h2aa == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28377); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28379 = 12'h2ab == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28378); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28380 = 12'h2ac == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28379); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28381 = 12'h2ad == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28380); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28382 = 12'h2ae == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28381); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28383 = 12'h2af == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28382); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28384 = 12'h2b0 == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28383); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28385 = 12'h2b1 == _T_837 ? $signed(-7'sh6) : $signed(_GEN_28384); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28386 = 12'h2b2 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28385); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28387 = 12'h2b3 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28386); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28388 = 12'h2b4 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28387); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28389 = 12'h2b5 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28388); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28390 = 12'h2b6 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28389); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28391 = 12'h2b7 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28390); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28392 = 12'h2b8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28391); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28393 = 12'h2b9 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28392); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28394 = 12'h2ba == _T_837 ? $signed(7'sh15) : $signed(_GEN_28393); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28395 = 12'h2bb == _T_837 ? $signed(7'sh14) : $signed(_GEN_28394); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28396 = 12'h2bc == _T_837 ? $signed(7'sh14) : $signed(_GEN_28395); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28397 = 12'h2bd == _T_837 ? $signed(7'sh13) : $signed(_GEN_28396); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28398 = 12'h2be == _T_837 ? $signed(7'sh12) : $signed(_GEN_28397); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28399 = 12'h2bf == _T_837 ? $signed(7'sh11) : $signed(_GEN_28398); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28400 = 12'h2c0 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28399); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28401 = 12'h2c1 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28400); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28402 = 12'h2c2 == _T_837 ? $signed(7'shf) : $signed(_GEN_28401); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28403 = 12'h2c3 == _T_837 ? $signed(7'shf) : $signed(_GEN_28402); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28404 = 12'h2c4 == _T_837 ? $signed(7'she) : $signed(_GEN_28403); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28405 = 12'h2c5 == _T_837 ? $signed(7'shd) : $signed(_GEN_28404); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28406 = 12'h2c6 == _T_837 ? $signed(7'shc) : $signed(_GEN_28405); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28407 = 12'h2c7 == _T_837 ? $signed(7'shc) : $signed(_GEN_28406); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28408 = 12'h2c8 == _T_837 ? $signed(7'shb) : $signed(_GEN_28407); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28409 = 12'h2c9 == _T_837 ? $signed(7'sha) : $signed(_GEN_28408); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28410 = 12'h2ca == _T_837 ? $signed(7'sha) : $signed(_GEN_28409); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28411 = 12'h2cb == _T_837 ? $signed(7'sh9) : $signed(_GEN_28410); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28412 = 12'h2cc == _T_837 ? $signed(7'sh8) : $signed(_GEN_28411); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28413 = 12'h2cd == _T_837 ? $signed(7'sh8) : $signed(_GEN_28412); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28414 = 12'h2ce == _T_837 ? $signed(7'sh7) : $signed(_GEN_28413); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28415 = 12'h2cf == _T_837 ? $signed(7'sh6) : $signed(_GEN_28414); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28416 = 12'h2d0 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28415); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28417 = 12'h2d1 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28416); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28418 = 12'h2d2 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28417); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28419 = 12'h2d3 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28418); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28420 = 12'h2d4 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28419); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28421 = 12'h2d5 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28420); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28422 = 12'h2d6 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28421); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28423 = 12'h2d7 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28422); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28424 = 12'h2d8 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28423); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28425 = 12'h2d9 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28424); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28426 = 12'h2da == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28425); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28427 = 12'h2db == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28426); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28428 = 12'h2dc == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28427); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28429 = 12'h2dd == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28428); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28430 = 12'h2de == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28429); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28431 = 12'h2df == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28430); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28432 = 12'h2e0 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28431); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28433 = 12'h2e1 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28432); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28434 = 12'h2e2 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28433); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28435 = 12'h2e3 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28434); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28436 = 12'h2e4 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28435); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28437 = 12'h2e5 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28436); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28438 = 12'h2e6 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28437); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28439 = 12'h2e7 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28438); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28440 = 12'h2e8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28439); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28441 = 12'h2e9 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28440); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28442 = 12'h2ea == _T_837 ? $signed(7'sh14) : $signed(_GEN_28441); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28443 = 12'h2eb == _T_837 ? $signed(7'sh14) : $signed(_GEN_28442); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28444 = 12'h2ec == _T_837 ? $signed(7'sh13) : $signed(_GEN_28443); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28445 = 12'h2ed == _T_837 ? $signed(7'sh12) : $signed(_GEN_28444); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28446 = 12'h2ee == _T_837 ? $signed(7'sh11) : $signed(_GEN_28445); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28447 = 12'h2ef == _T_837 ? $signed(7'sh11) : $signed(_GEN_28446); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28448 = 12'h2f0 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28447); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28449 = 12'h2f1 == _T_837 ? $signed(7'shf) : $signed(_GEN_28448); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28450 = 12'h2f2 == _T_837 ? $signed(7'shf) : $signed(_GEN_28449); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28451 = 12'h2f3 == _T_837 ? $signed(7'she) : $signed(_GEN_28450); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28452 = 12'h2f4 == _T_837 ? $signed(7'shd) : $signed(_GEN_28451); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28453 = 12'h2f5 == _T_837 ? $signed(7'shc) : $signed(_GEN_28452); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28454 = 12'h2f6 == _T_837 ? $signed(7'shc) : $signed(_GEN_28453); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28455 = 12'h2f7 == _T_837 ? $signed(7'shb) : $signed(_GEN_28454); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28456 = 12'h2f8 == _T_837 ? $signed(7'sha) : $signed(_GEN_28455); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28457 = 12'h2f9 == _T_837 ? $signed(7'sha) : $signed(_GEN_28456); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28458 = 12'h2fa == _T_837 ? $signed(7'sh9) : $signed(_GEN_28457); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28459 = 12'h2fb == _T_837 ? $signed(7'sh8) : $signed(_GEN_28458); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28460 = 12'h2fc == _T_837 ? $signed(7'sh8) : $signed(_GEN_28459); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28461 = 12'h2fd == _T_837 ? $signed(7'sh7) : $signed(_GEN_28460); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28462 = 12'h2fe == _T_837 ? $signed(7'sh6) : $signed(_GEN_28461); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28463 = 12'h2ff == _T_837 ? $signed(7'sh5) : $signed(_GEN_28462); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28464 = 12'h300 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28463); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28465 = 12'h301 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28464); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28466 = 12'h302 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28465); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28467 = 12'h303 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28466); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28468 = 12'h304 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28467); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28469 = 12'h305 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28468); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28470 = 12'h306 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28469); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28471 = 12'h307 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28470); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28472 = 12'h308 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28471); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28473 = 12'h309 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28472); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28474 = 12'h30a == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28473); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28475 = 12'h30b == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28474); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28476 = 12'h30c == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28475); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28477 = 12'h30d == _T_837 ? $signed(-7'sh5) : $signed(_GEN_28476); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28478 = 12'h30e == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28477); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28479 = 12'h30f == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28478); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28480 = 12'h310 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28479); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28481 = 12'h311 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28480); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28482 = 12'h312 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28481); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28483 = 12'h313 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28482); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28484 = 12'h314 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28483); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28485 = 12'h315 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28484); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28486 = 12'h316 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28485); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28487 = 12'h317 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28486); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28488 = 12'h318 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28487); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28489 = 12'h319 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28488); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28490 = 12'h31a == _T_837 ? $signed(7'sh14) : $signed(_GEN_28489); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28491 = 12'h31b == _T_837 ? $signed(7'sh13) : $signed(_GEN_28490); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28492 = 12'h31c == _T_837 ? $signed(7'sh12) : $signed(_GEN_28491); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28493 = 12'h31d == _T_837 ? $signed(7'sh11) : $signed(_GEN_28492); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28494 = 12'h31e == _T_837 ? $signed(7'sh11) : $signed(_GEN_28493); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28495 = 12'h31f == _T_837 ? $signed(7'sh10) : $signed(_GEN_28494); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28496 = 12'h320 == _T_837 ? $signed(7'shf) : $signed(_GEN_28495); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28497 = 12'h321 == _T_837 ? $signed(7'shf) : $signed(_GEN_28496); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28498 = 12'h322 == _T_837 ? $signed(7'she) : $signed(_GEN_28497); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28499 = 12'h323 == _T_837 ? $signed(7'shd) : $signed(_GEN_28498); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28500 = 12'h324 == _T_837 ? $signed(7'shc) : $signed(_GEN_28499); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28501 = 12'h325 == _T_837 ? $signed(7'shc) : $signed(_GEN_28500); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28502 = 12'h326 == _T_837 ? $signed(7'shb) : $signed(_GEN_28501); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28503 = 12'h327 == _T_837 ? $signed(7'sha) : $signed(_GEN_28502); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28504 = 12'h328 == _T_837 ? $signed(7'sha) : $signed(_GEN_28503); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28505 = 12'h329 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28504); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28506 = 12'h32a == _T_837 ? $signed(7'sh8) : $signed(_GEN_28505); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28507 = 12'h32b == _T_837 ? $signed(7'sh8) : $signed(_GEN_28506); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28508 = 12'h32c == _T_837 ? $signed(7'sh7) : $signed(_GEN_28507); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28509 = 12'h32d == _T_837 ? $signed(7'sh6) : $signed(_GEN_28508); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28510 = 12'h32e == _T_837 ? $signed(7'sh5) : $signed(_GEN_28509); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28511 = 12'h32f == _T_837 ? $signed(7'sh5) : $signed(_GEN_28510); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28512 = 12'h330 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28511); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28513 = 12'h331 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28512); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28514 = 12'h332 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28513); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28515 = 12'h333 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28514); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28516 = 12'h334 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28515); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28517 = 12'h335 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28516); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28518 = 12'h336 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28517); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28519 = 12'h337 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28518); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28520 = 12'h338 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28519); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28521 = 12'h339 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28520); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28522 = 12'h33a == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28521); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28523 = 12'h33b == _T_837 ? $signed(-7'sh4) : $signed(_GEN_28522); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28524 = 12'h33c == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28523); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28525 = 12'h33d == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28524); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28526 = 12'h33e == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28525); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28527 = 12'h33f == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28526); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28528 = 12'h340 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28527); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28529 = 12'h341 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28528); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28530 = 12'h342 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28529); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28531 = 12'h343 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28530); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28532 = 12'h344 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28531); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28533 = 12'h345 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28532); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28534 = 12'h346 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28533); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28535 = 12'h347 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28534); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28536 = 12'h348 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28535); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28537 = 12'h349 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28536); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28538 = 12'h34a == _T_837 ? $signed(7'sh13) : $signed(_GEN_28537); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28539 = 12'h34b == _T_837 ? $signed(7'sh12) : $signed(_GEN_28538); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28540 = 12'h34c == _T_837 ? $signed(7'sh11) : $signed(_GEN_28539); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28541 = 12'h34d == _T_837 ? $signed(7'sh11) : $signed(_GEN_28540); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28542 = 12'h34e == _T_837 ? $signed(7'sh10) : $signed(_GEN_28541); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28543 = 12'h34f == _T_837 ? $signed(7'shf) : $signed(_GEN_28542); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28544 = 12'h350 == _T_837 ? $signed(7'shf) : $signed(_GEN_28543); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28545 = 12'h351 == _T_837 ? $signed(7'she) : $signed(_GEN_28544); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28546 = 12'h352 == _T_837 ? $signed(7'shd) : $signed(_GEN_28545); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28547 = 12'h353 == _T_837 ? $signed(7'shc) : $signed(_GEN_28546); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28548 = 12'h354 == _T_837 ? $signed(7'shc) : $signed(_GEN_28547); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28549 = 12'h355 == _T_837 ? $signed(7'shb) : $signed(_GEN_28548); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28550 = 12'h356 == _T_837 ? $signed(7'sha) : $signed(_GEN_28549); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28551 = 12'h357 == _T_837 ? $signed(7'sha) : $signed(_GEN_28550); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28552 = 12'h358 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28551); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28553 = 12'h359 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28552); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28554 = 12'h35a == _T_837 ? $signed(7'sh8) : $signed(_GEN_28553); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28555 = 12'h35b == _T_837 ? $signed(7'sh7) : $signed(_GEN_28554); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28556 = 12'h35c == _T_837 ? $signed(7'sh6) : $signed(_GEN_28555); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28557 = 12'h35d == _T_837 ? $signed(7'sh5) : $signed(_GEN_28556); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28558 = 12'h35e == _T_837 ? $signed(7'sh5) : $signed(_GEN_28557); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28559 = 12'h35f == _T_837 ? $signed(7'sh4) : $signed(_GEN_28558); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28560 = 12'h360 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28559); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28561 = 12'h361 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28560); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28562 = 12'h362 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28561); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28563 = 12'h363 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28562); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28564 = 12'h364 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28563); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28565 = 12'h365 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28564); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28566 = 12'h366 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28565); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28567 = 12'h367 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28566); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28568 = 12'h368 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28567); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28569 = 12'h369 == _T_837 ? $signed(-7'sh3) : $signed(_GEN_28568); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28570 = 12'h36a == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28569); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28571 = 12'h36b == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28570); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28572 = 12'h36c == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28571); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28573 = 12'h36d == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28572); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28574 = 12'h36e == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28573); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28575 = 12'h36f == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28574); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28576 = 12'h370 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28575); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28577 = 12'h371 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28576); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28578 = 12'h372 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28577); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28579 = 12'h373 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28578); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28580 = 12'h374 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28579); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28581 = 12'h375 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28580); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28582 = 12'h376 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28581); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28583 = 12'h377 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28582); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28584 = 12'h378 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28583); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28585 = 12'h379 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28584); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28586 = 12'h37a == _T_837 ? $signed(7'sh12) : $signed(_GEN_28585); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28587 = 12'h37b == _T_837 ? $signed(7'sh11) : $signed(_GEN_28586); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28588 = 12'h37c == _T_837 ? $signed(7'sh11) : $signed(_GEN_28587); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28589 = 12'h37d == _T_837 ? $signed(7'sh10) : $signed(_GEN_28588); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28590 = 12'h37e == _T_837 ? $signed(7'shf) : $signed(_GEN_28589); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28591 = 12'h37f == _T_837 ? $signed(7'shf) : $signed(_GEN_28590); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28592 = 12'h380 == _T_837 ? $signed(7'she) : $signed(_GEN_28591); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28593 = 12'h381 == _T_837 ? $signed(7'shd) : $signed(_GEN_28592); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28594 = 12'h382 == _T_837 ? $signed(7'shc) : $signed(_GEN_28593); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28595 = 12'h383 == _T_837 ? $signed(7'shc) : $signed(_GEN_28594); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28596 = 12'h384 == _T_837 ? $signed(7'shb) : $signed(_GEN_28595); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28597 = 12'h385 == _T_837 ? $signed(7'sha) : $signed(_GEN_28596); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28598 = 12'h386 == _T_837 ? $signed(7'sha) : $signed(_GEN_28597); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28599 = 12'h387 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28598); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28600 = 12'h388 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28599); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28601 = 12'h389 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28600); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28602 = 12'h38a == _T_837 ? $signed(7'sh7) : $signed(_GEN_28601); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28603 = 12'h38b == _T_837 ? $signed(7'sh6) : $signed(_GEN_28602); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28604 = 12'h38c == _T_837 ? $signed(7'sh5) : $signed(_GEN_28603); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28605 = 12'h38d == _T_837 ? $signed(7'sh5) : $signed(_GEN_28604); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28606 = 12'h38e == _T_837 ? $signed(7'sh4) : $signed(_GEN_28605); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28607 = 12'h38f == _T_837 ? $signed(7'sh3) : $signed(_GEN_28606); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28608 = 12'h390 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28607); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28609 = 12'h391 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28608); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28610 = 12'h392 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28609); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28611 = 12'h393 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28610); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28612 = 12'h394 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28611); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28613 = 12'h395 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28612); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28614 = 12'h396 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28613); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28615 = 12'h397 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28614); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28616 = 12'h398 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28615); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28617 = 12'h399 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28616); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28618 = 12'h39a == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28617); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28619 = 12'h39b == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28618); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28620 = 12'h39c == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28619); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28621 = 12'h39d == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28620); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28622 = 12'h39e == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28621); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28623 = 12'h39f == _T_837 ? $signed(7'sh19) : $signed(_GEN_28622); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28624 = 12'h3a0 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28623); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28625 = 12'h3a1 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28624); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28626 = 12'h3a2 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28625); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28627 = 12'h3a3 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28626); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28628 = 12'h3a4 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28627); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28629 = 12'h3a5 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28628); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28630 = 12'h3a6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28629); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28631 = 12'h3a7 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28630); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28632 = 12'h3a8 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28631); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28633 = 12'h3a9 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28632); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28634 = 12'h3aa == _T_837 ? $signed(7'sh11) : $signed(_GEN_28633); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28635 = 12'h3ab == _T_837 ? $signed(7'sh11) : $signed(_GEN_28634); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28636 = 12'h3ac == _T_837 ? $signed(7'sh10) : $signed(_GEN_28635); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28637 = 12'h3ad == _T_837 ? $signed(7'shf) : $signed(_GEN_28636); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28638 = 12'h3ae == _T_837 ? $signed(7'shf) : $signed(_GEN_28637); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28639 = 12'h3af == _T_837 ? $signed(7'she) : $signed(_GEN_28638); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28640 = 12'h3b0 == _T_837 ? $signed(7'shd) : $signed(_GEN_28639); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28641 = 12'h3b1 == _T_837 ? $signed(7'shc) : $signed(_GEN_28640); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28642 = 12'h3b2 == _T_837 ? $signed(7'shc) : $signed(_GEN_28641); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28643 = 12'h3b3 == _T_837 ? $signed(7'shb) : $signed(_GEN_28642); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28644 = 12'h3b4 == _T_837 ? $signed(7'sha) : $signed(_GEN_28643); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28645 = 12'h3b5 == _T_837 ? $signed(7'sha) : $signed(_GEN_28644); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28646 = 12'h3b6 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28645); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28647 = 12'h3b7 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28646); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28648 = 12'h3b8 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28647); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28649 = 12'h3b9 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28648); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28650 = 12'h3ba == _T_837 ? $signed(7'sh6) : $signed(_GEN_28649); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28651 = 12'h3bb == _T_837 ? $signed(7'sh5) : $signed(_GEN_28650); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28652 = 12'h3bc == _T_837 ? $signed(7'sh5) : $signed(_GEN_28651); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28653 = 12'h3bd == _T_837 ? $signed(7'sh4) : $signed(_GEN_28652); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28654 = 12'h3be == _T_837 ? $signed(7'sh3) : $signed(_GEN_28653); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28655 = 12'h3bf == _T_837 ? $signed(7'sh3) : $signed(_GEN_28654); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28656 = 12'h3c0 == _T_837 ? $signed(7'sh2) : $signed(_GEN_28655); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28657 = 12'h3c1 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28656); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28658 = 12'h3c2 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28657); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28659 = 12'h3c3 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28658); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28660 = 12'h3c4 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28659); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28661 = 12'h3c5 == _T_837 ? $signed(-7'sh2) : $signed(_GEN_28660); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28662 = 12'h3c6 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28661); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28663 = 12'h3c7 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28662); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28664 = 12'h3c8 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28663); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28665 = 12'h3c9 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28664); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28666 = 12'h3ca == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28665); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28667 = 12'h3cb == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28666); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28668 = 12'h3cc == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28667); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28669 = 12'h3cd == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28668); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28670 = 12'h3ce == _T_837 ? $signed(7'sh19) : $signed(_GEN_28669); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28671 = 12'h3cf == _T_837 ? $signed(7'sh18) : $signed(_GEN_28670); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28672 = 12'h3d0 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28671); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28673 = 12'h3d1 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28672); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28674 = 12'h3d2 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28673); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28675 = 12'h3d3 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28674); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28676 = 12'h3d4 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28675); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28677 = 12'h3d5 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28676); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28678 = 12'h3d6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28677); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28679 = 12'h3d7 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28678); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28680 = 12'h3d8 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28679); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28681 = 12'h3d9 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28680); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28682 = 12'h3da == _T_837 ? $signed(7'sh11) : $signed(_GEN_28681); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28683 = 12'h3db == _T_837 ? $signed(7'sh10) : $signed(_GEN_28682); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28684 = 12'h3dc == _T_837 ? $signed(7'shf) : $signed(_GEN_28683); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28685 = 12'h3dd == _T_837 ? $signed(7'shf) : $signed(_GEN_28684); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28686 = 12'h3de == _T_837 ? $signed(7'she) : $signed(_GEN_28685); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28687 = 12'h3df == _T_837 ? $signed(7'shd) : $signed(_GEN_28686); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28688 = 12'h3e0 == _T_837 ? $signed(7'shc) : $signed(_GEN_28687); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28689 = 12'h3e1 == _T_837 ? $signed(7'shc) : $signed(_GEN_28688); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28690 = 12'h3e2 == _T_837 ? $signed(7'shb) : $signed(_GEN_28689); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28691 = 12'h3e3 == _T_837 ? $signed(7'sha) : $signed(_GEN_28690); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28692 = 12'h3e4 == _T_837 ? $signed(7'sha) : $signed(_GEN_28691); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28693 = 12'h3e5 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28692); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28694 = 12'h3e6 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28693); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28695 = 12'h3e7 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28694); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28696 = 12'h3e8 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28695); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28697 = 12'h3e9 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28696); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28698 = 12'h3ea == _T_837 ? $signed(7'sh5) : $signed(_GEN_28697); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28699 = 12'h3eb == _T_837 ? $signed(7'sh5) : $signed(_GEN_28698); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28700 = 12'h3ec == _T_837 ? $signed(7'sh4) : $signed(_GEN_28699); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28701 = 12'h3ed == _T_837 ? $signed(7'sh3) : $signed(_GEN_28700); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28702 = 12'h3ee == _T_837 ? $signed(7'sh3) : $signed(_GEN_28701); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28703 = 12'h3ef == _T_837 ? $signed(7'sh2) : $signed(_GEN_28702); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28704 = 12'h3f0 == _T_837 ? $signed(7'sh1) : $signed(_GEN_28703); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28705 = 12'h3f1 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28704); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28706 = 12'h3f2 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28705); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28707 = 12'h3f3 == _T_837 ? $signed(-7'sh1) : $signed(_GEN_28706); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28708 = 12'h3f4 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28707); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28709 = 12'h3f5 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28708); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28710 = 12'h3f6 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28709); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28711 = 12'h3f7 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28710); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28712 = 12'h3f8 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28711); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28713 = 12'h3f9 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28712); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28714 = 12'h3fa == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28713); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28715 = 12'h3fb == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28714); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28716 = 12'h3fc == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28715); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28717 = 12'h3fd == _T_837 ? $signed(7'sh19) : $signed(_GEN_28716); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28718 = 12'h3fe == _T_837 ? $signed(7'sh18) : $signed(_GEN_28717); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28719 = 12'h3ff == _T_837 ? $signed(7'sh18) : $signed(_GEN_28718); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28720 = 12'h400 == _T_837 ? $signed(7'sh17) : $signed(_GEN_28719); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28721 = 12'h401 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28720); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28722 = 12'h402 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28721); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28723 = 12'h403 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28722); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28724 = 12'h404 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28723); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28725 = 12'h405 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28724); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28726 = 12'h406 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28725); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28727 = 12'h407 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28726); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28728 = 12'h408 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28727); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28729 = 12'h409 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28728); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28730 = 12'h40a == _T_837 ? $signed(7'sh10) : $signed(_GEN_28729); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28731 = 12'h40b == _T_837 ? $signed(7'shf) : $signed(_GEN_28730); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28732 = 12'h40c == _T_837 ? $signed(7'shf) : $signed(_GEN_28731); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28733 = 12'h40d == _T_837 ? $signed(7'she) : $signed(_GEN_28732); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28734 = 12'h40e == _T_837 ? $signed(7'shd) : $signed(_GEN_28733); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28735 = 12'h40f == _T_837 ? $signed(7'shc) : $signed(_GEN_28734); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28736 = 12'h410 == _T_837 ? $signed(7'shc) : $signed(_GEN_28735); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28737 = 12'h411 == _T_837 ? $signed(7'shb) : $signed(_GEN_28736); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28738 = 12'h412 == _T_837 ? $signed(7'sha) : $signed(_GEN_28737); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28739 = 12'h413 == _T_837 ? $signed(7'sha) : $signed(_GEN_28738); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28740 = 12'h414 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28739); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28741 = 12'h415 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28740); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28742 = 12'h416 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28741); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28743 = 12'h417 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28742); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28744 = 12'h418 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28743); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28745 = 12'h419 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28744); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28746 = 12'h41a == _T_837 ? $signed(7'sh5) : $signed(_GEN_28745); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28747 = 12'h41b == _T_837 ? $signed(7'sh4) : $signed(_GEN_28746); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28748 = 12'h41c == _T_837 ? $signed(7'sh3) : $signed(_GEN_28747); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28749 = 12'h41d == _T_837 ? $signed(7'sh3) : $signed(_GEN_28748); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28750 = 12'h41e == _T_837 ? $signed(7'sh2) : $signed(_GEN_28749); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28751 = 12'h41f == _T_837 ? $signed(7'sh1) : $signed(_GEN_28750); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28752 = 12'h420 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28751); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28753 = 12'h421 == _T_837 ? $signed(7'sh0) : $signed(_GEN_28752); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28754 = 12'h422 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28753); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28755 = 12'h423 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28754); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28756 = 12'h424 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28755); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28757 = 12'h425 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28756); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28758 = 12'h426 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28757); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28759 = 12'h427 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28758); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28760 = 12'h428 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28759); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28761 = 12'h429 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28760); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28762 = 12'h42a == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28761); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28763 = 12'h42b == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28762); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28764 = 12'h42c == _T_837 ? $signed(7'sh19) : $signed(_GEN_28763); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28765 = 12'h42d == _T_837 ? $signed(7'sh18) : $signed(_GEN_28764); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28766 = 12'h42e == _T_837 ? $signed(7'sh18) : $signed(_GEN_28765); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28767 = 12'h42f == _T_837 ? $signed(7'sh17) : $signed(_GEN_28766); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28768 = 12'h430 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28767); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28769 = 12'h431 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28768); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28770 = 12'h432 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28769); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28771 = 12'h433 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28770); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28772 = 12'h434 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28771); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28773 = 12'h435 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28772); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28774 = 12'h436 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28773); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28775 = 12'h437 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28774); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28776 = 12'h438 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28775); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28777 = 12'h439 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28776); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28778 = 12'h43a == _T_837 ? $signed(7'shf) : $signed(_GEN_28777); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28779 = 12'h43b == _T_837 ? $signed(7'shf) : $signed(_GEN_28778); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28780 = 12'h43c == _T_837 ? $signed(7'she) : $signed(_GEN_28779); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28781 = 12'h43d == _T_837 ? $signed(7'shd) : $signed(_GEN_28780); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28782 = 12'h43e == _T_837 ? $signed(7'shc) : $signed(_GEN_28781); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28783 = 12'h43f == _T_837 ? $signed(7'shc) : $signed(_GEN_28782); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28784 = 12'h440 == _T_837 ? $signed(7'shb) : $signed(_GEN_28783); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28785 = 12'h441 == _T_837 ? $signed(7'sha) : $signed(_GEN_28784); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28786 = 12'h442 == _T_837 ? $signed(7'sha) : $signed(_GEN_28785); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28787 = 12'h443 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28786); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28788 = 12'h444 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28787); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28789 = 12'h445 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28788); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28790 = 12'h446 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28789); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28791 = 12'h447 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28790); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28792 = 12'h448 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28791); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28793 = 12'h449 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28792); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28794 = 12'h44a == _T_837 ? $signed(7'sh4) : $signed(_GEN_28793); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28795 = 12'h44b == _T_837 ? $signed(7'sh3) : $signed(_GEN_28794); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28796 = 12'h44c == _T_837 ? $signed(7'sh3) : $signed(_GEN_28795); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28797 = 12'h44d == _T_837 ? $signed(7'sh2) : $signed(_GEN_28796); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28798 = 12'h44e == _T_837 ? $signed(7'sh1) : $signed(_GEN_28797); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28799 = 12'h44f == _T_837 ? $signed(7'sh0) : $signed(_GEN_28798); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28800 = 12'h450 == _T_837 ? $signed(7'sh21) : $signed(_GEN_28799); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28801 = 12'h451 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28800); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28802 = 12'h452 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28801); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28803 = 12'h453 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28802); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28804 = 12'h454 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28803); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28805 = 12'h455 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28804); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28806 = 12'h456 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28805); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28807 = 12'h457 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28806); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28808 = 12'h458 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28807); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28809 = 12'h459 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28808); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28810 = 12'h45a == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28809); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28811 = 12'h45b == _T_837 ? $signed(7'sh19) : $signed(_GEN_28810); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28812 = 12'h45c == _T_837 ? $signed(7'sh18) : $signed(_GEN_28811); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28813 = 12'h45d == _T_837 ? $signed(7'sh18) : $signed(_GEN_28812); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28814 = 12'h45e == _T_837 ? $signed(7'sh17) : $signed(_GEN_28813); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28815 = 12'h45f == _T_837 ? $signed(7'sh16) : $signed(_GEN_28814); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28816 = 12'h460 == _T_837 ? $signed(7'sh16) : $signed(_GEN_28815); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28817 = 12'h461 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28816); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28818 = 12'h462 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28817); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28819 = 12'h463 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28818); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28820 = 12'h464 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28819); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28821 = 12'h465 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28820); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28822 = 12'h466 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28821); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28823 = 12'h467 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28822); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28824 = 12'h468 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28823); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28825 = 12'h469 == _T_837 ? $signed(7'shf) : $signed(_GEN_28824); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28826 = 12'h46a == _T_837 ? $signed(7'shf) : $signed(_GEN_28825); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28827 = 12'h46b == _T_837 ? $signed(7'she) : $signed(_GEN_28826); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28828 = 12'h46c == _T_837 ? $signed(7'shd) : $signed(_GEN_28827); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28829 = 12'h46d == _T_837 ? $signed(7'shc) : $signed(_GEN_28828); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28830 = 12'h46e == _T_837 ? $signed(7'shc) : $signed(_GEN_28829); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28831 = 12'h46f == _T_837 ? $signed(7'shb) : $signed(_GEN_28830); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28832 = 12'h470 == _T_837 ? $signed(7'sha) : $signed(_GEN_28831); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28833 = 12'h471 == _T_837 ? $signed(7'sha) : $signed(_GEN_28832); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28834 = 12'h472 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28833); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28835 = 12'h473 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28834); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28836 = 12'h474 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28835); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28837 = 12'h475 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28836); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28838 = 12'h476 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28837); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28839 = 12'h477 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28838); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28840 = 12'h478 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28839); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28841 = 12'h479 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28840); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28842 = 12'h47a == _T_837 ? $signed(7'sh3) : $signed(_GEN_28841); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28843 = 12'h47b == _T_837 ? $signed(7'sh3) : $signed(_GEN_28842); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28844 = 12'h47c == _T_837 ? $signed(7'sh2) : $signed(_GEN_28843); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28845 = 12'h47d == _T_837 ? $signed(7'sh1) : $signed(_GEN_28844); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28846 = 12'h47e == _T_837 ? $signed(7'sh22) : $signed(_GEN_28845); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28847 = 12'h47f == _T_837 ? $signed(7'sh21) : $signed(_GEN_28846); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28848 = 12'h480 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28847); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28849 = 12'h481 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28848); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28850 = 12'h482 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28849); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28851 = 12'h483 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28850); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28852 = 12'h484 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28851); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28853 = 12'h485 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28852); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28854 = 12'h486 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28853); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28855 = 12'h487 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28854); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28856 = 12'h488 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28855); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28857 = 12'h489 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28856); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28858 = 12'h48a == _T_837 ? $signed(7'sh19) : $signed(_GEN_28857); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28859 = 12'h48b == _T_837 ? $signed(7'sh18) : $signed(_GEN_28858); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28860 = 12'h48c == _T_837 ? $signed(7'sh18) : $signed(_GEN_28859); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28861 = 12'h48d == _T_837 ? $signed(7'sh17) : $signed(_GEN_28860); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28862 = 12'h48e == _T_837 ? $signed(7'sh16) : $signed(_GEN_28861); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28863 = 12'h48f == _T_837 ? $signed(7'sh16) : $signed(_GEN_28862); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28864 = 12'h490 == _T_837 ? $signed(7'sh15) : $signed(_GEN_28863); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28865 = 12'h491 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28864); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28866 = 12'h492 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28865); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28867 = 12'h493 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28866); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28868 = 12'h494 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28867); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28869 = 12'h495 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28868); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28870 = 12'h496 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28869); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28871 = 12'h497 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28870); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28872 = 12'h498 == _T_837 ? $signed(7'shf) : $signed(_GEN_28871); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28873 = 12'h499 == _T_837 ? $signed(7'shf) : $signed(_GEN_28872); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28874 = 12'h49a == _T_837 ? $signed(7'she) : $signed(_GEN_28873); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28875 = 12'h49b == _T_837 ? $signed(7'shd) : $signed(_GEN_28874); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28876 = 12'h49c == _T_837 ? $signed(7'shc) : $signed(_GEN_28875); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28877 = 12'h49d == _T_837 ? $signed(7'shc) : $signed(_GEN_28876); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28878 = 12'h49e == _T_837 ? $signed(7'shb) : $signed(_GEN_28877); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28879 = 12'h49f == _T_837 ? $signed(7'sha) : $signed(_GEN_28878); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28880 = 12'h4a0 == _T_837 ? $signed(7'sha) : $signed(_GEN_28879); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28881 = 12'h4a1 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28880); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28882 = 12'h4a2 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28881); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28883 = 12'h4a3 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28882); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28884 = 12'h4a4 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28883); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28885 = 12'h4a5 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28884); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28886 = 12'h4a6 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28885); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28887 = 12'h4a7 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28886); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28888 = 12'h4a8 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28887); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28889 = 12'h4a9 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28888); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28890 = 12'h4aa == _T_837 ? $signed(7'sh3) : $signed(_GEN_28889); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28891 = 12'h4ab == _T_837 ? $signed(7'sh2) : $signed(_GEN_28890); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28892 = 12'h4ac == _T_837 ? $signed(7'sh22) : $signed(_GEN_28891); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28893 = 12'h4ad == _T_837 ? $signed(7'sh22) : $signed(_GEN_28892); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28894 = 12'h4ae == _T_837 ? $signed(7'sh21) : $signed(_GEN_28893); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28895 = 12'h4af == _T_837 ? $signed(7'sh20) : $signed(_GEN_28894); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28896 = 12'h4b0 == _T_837 ? $signed(7'sh20) : $signed(_GEN_28895); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28897 = 12'h4b1 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28896); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28898 = 12'h4b2 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28897); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28899 = 12'h4b3 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28898); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28900 = 12'h4b4 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28899); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28901 = 12'h4b5 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28900); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28902 = 12'h4b6 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28901); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28903 = 12'h4b7 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28902); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28904 = 12'h4b8 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28903); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28905 = 12'h4b9 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28904); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28906 = 12'h4ba == _T_837 ? $signed(7'sh18) : $signed(_GEN_28905); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28907 = 12'h4bb == _T_837 ? $signed(7'sh18) : $signed(_GEN_28906); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28908 = 12'h4bc == _T_837 ? $signed(7'sh17) : $signed(_GEN_28907); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28909 = 12'h4bd == _T_837 ? $signed(7'sh16) : $signed(_GEN_28908); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28910 = 12'h4be == _T_837 ? $signed(7'sh16) : $signed(_GEN_28909); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28911 = 12'h4bf == _T_837 ? $signed(7'sh15) : $signed(_GEN_28910); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28912 = 12'h4c0 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28911); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28913 = 12'h4c1 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28912); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28914 = 12'h4c2 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28913); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28915 = 12'h4c3 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28914); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28916 = 12'h4c4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28915); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28917 = 12'h4c5 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28916); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28918 = 12'h4c6 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28917); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28919 = 12'h4c7 == _T_837 ? $signed(7'shf) : $signed(_GEN_28918); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28920 = 12'h4c8 == _T_837 ? $signed(7'shf) : $signed(_GEN_28919); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28921 = 12'h4c9 == _T_837 ? $signed(7'she) : $signed(_GEN_28920); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28922 = 12'h4ca == _T_837 ? $signed(7'shd) : $signed(_GEN_28921); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28923 = 12'h4cb == _T_837 ? $signed(7'shc) : $signed(_GEN_28922); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28924 = 12'h4cc == _T_837 ? $signed(7'shc) : $signed(_GEN_28923); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28925 = 12'h4cd == _T_837 ? $signed(7'shb) : $signed(_GEN_28924); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28926 = 12'h4ce == _T_837 ? $signed(7'sha) : $signed(_GEN_28925); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28927 = 12'h4cf == _T_837 ? $signed(7'sha) : $signed(_GEN_28926); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28928 = 12'h4d0 == _T_837 ? $signed(7'sh9) : $signed(_GEN_28927); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28929 = 12'h4d1 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28928); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28930 = 12'h4d2 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28929); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28931 = 12'h4d3 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28930); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28932 = 12'h4d4 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28931); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28933 = 12'h4d5 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28932); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28934 = 12'h4d6 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28933); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28935 = 12'h4d7 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28934); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28936 = 12'h4d8 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28935); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28937 = 12'h4d9 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28936); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28938 = 12'h4da == _T_837 ? $signed(7'sh23) : $signed(_GEN_28937); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28939 = 12'h4db == _T_837 ? $signed(7'sh22) : $signed(_GEN_28938); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28940 = 12'h4dc == _T_837 ? $signed(7'sh22) : $signed(_GEN_28939); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28941 = 12'h4dd == _T_837 ? $signed(7'sh21) : $signed(_GEN_28940); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28942 = 12'h4de == _T_837 ? $signed(7'sh20) : $signed(_GEN_28941); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28943 = 12'h4df == _T_837 ? $signed(7'sh20) : $signed(_GEN_28942); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28944 = 12'h4e0 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28943); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28945 = 12'h4e1 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28944); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28946 = 12'h4e2 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28945); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28947 = 12'h4e3 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28946); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28948 = 12'h4e4 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28947); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28949 = 12'h4e5 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28948); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28950 = 12'h4e6 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28949); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28951 = 12'h4e7 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28950); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28952 = 12'h4e8 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28951); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28953 = 12'h4e9 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28952); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28954 = 12'h4ea == _T_837 ? $signed(7'sh18) : $signed(_GEN_28953); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28955 = 12'h4eb == _T_837 ? $signed(7'sh17) : $signed(_GEN_28954); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28956 = 12'h4ec == _T_837 ? $signed(7'sh16) : $signed(_GEN_28955); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28957 = 12'h4ed == _T_837 ? $signed(7'sh16) : $signed(_GEN_28956); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28958 = 12'h4ee == _T_837 ? $signed(7'sh15) : $signed(_GEN_28957); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28959 = 12'h4ef == _T_837 ? $signed(7'sh14) : $signed(_GEN_28958); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28960 = 12'h4f0 == _T_837 ? $signed(7'sh14) : $signed(_GEN_28959); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28961 = 12'h4f1 == _T_837 ? $signed(7'sh13) : $signed(_GEN_28960); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28962 = 12'h4f2 == _T_837 ? $signed(7'sh12) : $signed(_GEN_28961); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28963 = 12'h4f3 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28962); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28964 = 12'h4f4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_28963); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28965 = 12'h4f5 == _T_837 ? $signed(7'sh10) : $signed(_GEN_28964); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28966 = 12'h4f6 == _T_837 ? $signed(7'shf) : $signed(_GEN_28965); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28967 = 12'h4f7 == _T_837 ? $signed(7'shf) : $signed(_GEN_28966); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28968 = 12'h4f8 == _T_837 ? $signed(7'she) : $signed(_GEN_28967); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28969 = 12'h4f9 == _T_837 ? $signed(7'shd) : $signed(_GEN_28968); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28970 = 12'h4fa == _T_837 ? $signed(7'shc) : $signed(_GEN_28969); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28971 = 12'h4fb == _T_837 ? $signed(7'shc) : $signed(_GEN_28970); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28972 = 12'h4fc == _T_837 ? $signed(7'shb) : $signed(_GEN_28971); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28973 = 12'h4fd == _T_837 ? $signed(7'sha) : $signed(_GEN_28972); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28974 = 12'h4fe == _T_837 ? $signed(7'sha) : $signed(_GEN_28973); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28975 = 12'h4ff == _T_837 ? $signed(7'sh9) : $signed(_GEN_28974); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28976 = 12'h500 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28975); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28977 = 12'h501 == _T_837 ? $signed(7'sh8) : $signed(_GEN_28976); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28978 = 12'h502 == _T_837 ? $signed(7'sh7) : $signed(_GEN_28977); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28979 = 12'h503 == _T_837 ? $signed(7'sh6) : $signed(_GEN_28978); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28980 = 12'h504 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28979); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28981 = 12'h505 == _T_837 ? $signed(7'sh5) : $signed(_GEN_28980); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28982 = 12'h506 == _T_837 ? $signed(7'sh4) : $signed(_GEN_28981); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28983 = 12'h507 == _T_837 ? $signed(7'sh3) : $signed(_GEN_28982); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28984 = 12'h508 == _T_837 ? $signed(7'sh24) : $signed(_GEN_28983); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28985 = 12'h509 == _T_837 ? $signed(7'sh23) : $signed(_GEN_28984); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28986 = 12'h50a == _T_837 ? $signed(7'sh22) : $signed(_GEN_28985); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28987 = 12'h50b == _T_837 ? $signed(7'sh22) : $signed(_GEN_28986); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28988 = 12'h50c == _T_837 ? $signed(7'sh21) : $signed(_GEN_28987); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28989 = 12'h50d == _T_837 ? $signed(7'sh20) : $signed(_GEN_28988); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28990 = 12'h50e == _T_837 ? $signed(7'sh20) : $signed(_GEN_28989); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28991 = 12'h50f == _T_837 ? $signed(7'sh1f) : $signed(_GEN_28990); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28992 = 12'h510 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_28991); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28993 = 12'h511 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28992); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28994 = 12'h512 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_28993); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28995 = 12'h513 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_28994); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28996 = 12'h514 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28995); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28997 = 12'h515 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_28996); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28998 = 12'h516 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_28997); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_28999 = 12'h517 == _T_837 ? $signed(7'sh19) : $signed(_GEN_28998); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29000 = 12'h518 == _T_837 ? $signed(7'sh18) : $signed(_GEN_28999); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29001 = 12'h519 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29000); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29002 = 12'h51a == _T_837 ? $signed(7'sh17) : $signed(_GEN_29001); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29003 = 12'h51b == _T_837 ? $signed(7'sh16) : $signed(_GEN_29002); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29004 = 12'h51c == _T_837 ? $signed(7'sh16) : $signed(_GEN_29003); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29005 = 12'h51d == _T_837 ? $signed(7'sh15) : $signed(_GEN_29004); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29006 = 12'h51e == _T_837 ? $signed(7'sh14) : $signed(_GEN_29005); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29007 = 12'h51f == _T_837 ? $signed(7'sh14) : $signed(_GEN_29006); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29008 = 12'h520 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29007); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29009 = 12'h521 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29008); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29010 = 12'h522 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29009); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29011 = 12'h523 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29010); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29012 = 12'h524 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29011); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29013 = 12'h525 == _T_837 ? $signed(7'shf) : $signed(_GEN_29012); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29014 = 12'h526 == _T_837 ? $signed(7'shf) : $signed(_GEN_29013); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29015 = 12'h527 == _T_837 ? $signed(7'she) : $signed(_GEN_29014); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29016 = 12'h528 == _T_837 ? $signed(7'shd) : $signed(_GEN_29015); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29017 = 12'h529 == _T_837 ? $signed(7'shc) : $signed(_GEN_29016); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29018 = 12'h52a == _T_837 ? $signed(7'shc) : $signed(_GEN_29017); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29019 = 12'h52b == _T_837 ? $signed(7'shb) : $signed(_GEN_29018); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29020 = 12'h52c == _T_837 ? $signed(7'sha) : $signed(_GEN_29019); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29021 = 12'h52d == _T_837 ? $signed(7'sha) : $signed(_GEN_29020); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29022 = 12'h52e == _T_837 ? $signed(7'sh9) : $signed(_GEN_29021); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29023 = 12'h52f == _T_837 ? $signed(7'sh8) : $signed(_GEN_29022); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29024 = 12'h530 == _T_837 ? $signed(7'sh8) : $signed(_GEN_29023); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29025 = 12'h531 == _T_837 ? $signed(7'sh7) : $signed(_GEN_29024); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29026 = 12'h532 == _T_837 ? $signed(7'sh6) : $signed(_GEN_29025); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29027 = 12'h533 == _T_837 ? $signed(7'sh5) : $signed(_GEN_29026); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29028 = 12'h534 == _T_837 ? $signed(7'sh5) : $signed(_GEN_29027); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29029 = 12'h535 == _T_837 ? $signed(7'sh4) : $signed(_GEN_29028); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29030 = 12'h536 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29029); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29031 = 12'h537 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29030); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29032 = 12'h538 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29031); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29033 = 12'h539 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29032); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29034 = 12'h53a == _T_837 ? $signed(7'sh22) : $signed(_GEN_29033); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29035 = 12'h53b == _T_837 ? $signed(7'sh21) : $signed(_GEN_29034); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29036 = 12'h53c == _T_837 ? $signed(7'sh20) : $signed(_GEN_29035); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29037 = 12'h53d == _T_837 ? $signed(7'sh20) : $signed(_GEN_29036); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29038 = 12'h53e == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29037); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29039 = 12'h53f == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29038); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29040 = 12'h540 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29039); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29041 = 12'h541 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29040); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29042 = 12'h542 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29041); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29043 = 12'h543 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29042); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29044 = 12'h544 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29043); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29045 = 12'h545 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29044); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29046 = 12'h546 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29045); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29047 = 12'h547 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29046); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29048 = 12'h548 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29047); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29049 = 12'h549 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29048); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29050 = 12'h54a == _T_837 ? $signed(7'sh16) : $signed(_GEN_29049); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29051 = 12'h54b == _T_837 ? $signed(7'sh16) : $signed(_GEN_29050); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29052 = 12'h54c == _T_837 ? $signed(7'sh15) : $signed(_GEN_29051); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29053 = 12'h54d == _T_837 ? $signed(7'sh14) : $signed(_GEN_29052); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29054 = 12'h54e == _T_837 ? $signed(7'sh14) : $signed(_GEN_29053); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29055 = 12'h54f == _T_837 ? $signed(7'sh13) : $signed(_GEN_29054); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29056 = 12'h550 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29055); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29057 = 12'h551 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29056); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29058 = 12'h552 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29057); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29059 = 12'h553 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29058); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29060 = 12'h554 == _T_837 ? $signed(7'shf) : $signed(_GEN_29059); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29061 = 12'h555 == _T_837 ? $signed(7'shf) : $signed(_GEN_29060); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29062 = 12'h556 == _T_837 ? $signed(7'she) : $signed(_GEN_29061); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29063 = 12'h557 == _T_837 ? $signed(7'shd) : $signed(_GEN_29062); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29064 = 12'h558 == _T_837 ? $signed(7'shc) : $signed(_GEN_29063); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29065 = 12'h559 == _T_837 ? $signed(7'shc) : $signed(_GEN_29064); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29066 = 12'h55a == _T_837 ? $signed(7'shb) : $signed(_GEN_29065); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29067 = 12'h55b == _T_837 ? $signed(7'sha) : $signed(_GEN_29066); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29068 = 12'h55c == _T_837 ? $signed(7'sha) : $signed(_GEN_29067); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29069 = 12'h55d == _T_837 ? $signed(7'sh9) : $signed(_GEN_29068); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29070 = 12'h55e == _T_837 ? $signed(7'sh8) : $signed(_GEN_29069); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29071 = 12'h55f == _T_837 ? $signed(7'sh8) : $signed(_GEN_29070); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29072 = 12'h560 == _T_837 ? $signed(7'sh7) : $signed(_GEN_29071); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29073 = 12'h561 == _T_837 ? $signed(7'sh6) : $signed(_GEN_29072); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29074 = 12'h562 == _T_837 ? $signed(7'sh5) : $signed(_GEN_29073); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29075 = 12'h563 == _T_837 ? $signed(7'sh5) : $signed(_GEN_29074); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29076 = 12'h564 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29075); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29077 = 12'h565 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29076); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29078 = 12'h566 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29077); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29079 = 12'h567 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29078); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29080 = 12'h568 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29079); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29081 = 12'h569 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29080); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29082 = 12'h56a == _T_837 ? $signed(7'sh21) : $signed(_GEN_29081); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29083 = 12'h56b == _T_837 ? $signed(7'sh20) : $signed(_GEN_29082); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29084 = 12'h56c == _T_837 ? $signed(7'sh20) : $signed(_GEN_29083); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29085 = 12'h56d == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29084); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29086 = 12'h56e == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29085); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29087 = 12'h56f == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29086); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29088 = 12'h570 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29087); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29089 = 12'h571 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29088); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29090 = 12'h572 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29089); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29091 = 12'h573 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29090); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29092 = 12'h574 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29091); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29093 = 12'h575 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29092); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29094 = 12'h576 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29093); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29095 = 12'h577 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29094); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29096 = 12'h578 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29095); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29097 = 12'h579 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29096); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29098 = 12'h57a == _T_837 ? $signed(7'sh16) : $signed(_GEN_29097); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29099 = 12'h57b == _T_837 ? $signed(7'sh15) : $signed(_GEN_29098); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29100 = 12'h57c == _T_837 ? $signed(7'sh14) : $signed(_GEN_29099); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29101 = 12'h57d == _T_837 ? $signed(7'sh14) : $signed(_GEN_29100); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29102 = 12'h57e == _T_837 ? $signed(7'sh13) : $signed(_GEN_29101); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29103 = 12'h57f == _T_837 ? $signed(7'sh12) : $signed(_GEN_29102); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29104 = 12'h580 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29103); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29105 = 12'h581 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29104); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29106 = 12'h582 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29105); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29107 = 12'h583 == _T_837 ? $signed(7'shf) : $signed(_GEN_29106); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29108 = 12'h584 == _T_837 ? $signed(7'shf) : $signed(_GEN_29107); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29109 = 12'h585 == _T_837 ? $signed(7'she) : $signed(_GEN_29108); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29110 = 12'h586 == _T_837 ? $signed(7'shd) : $signed(_GEN_29109); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29111 = 12'h587 == _T_837 ? $signed(7'shc) : $signed(_GEN_29110); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29112 = 12'h588 == _T_837 ? $signed(7'shc) : $signed(_GEN_29111); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29113 = 12'h589 == _T_837 ? $signed(7'shb) : $signed(_GEN_29112); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29114 = 12'h58a == _T_837 ? $signed(7'sha) : $signed(_GEN_29113); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29115 = 12'h58b == _T_837 ? $signed(7'sha) : $signed(_GEN_29114); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29116 = 12'h58c == _T_837 ? $signed(7'sh9) : $signed(_GEN_29115); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29117 = 12'h58d == _T_837 ? $signed(7'sh8) : $signed(_GEN_29116); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29118 = 12'h58e == _T_837 ? $signed(7'sh8) : $signed(_GEN_29117); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29119 = 12'h58f == _T_837 ? $signed(7'sh7) : $signed(_GEN_29118); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29120 = 12'h590 == _T_837 ? $signed(7'sh6) : $signed(_GEN_29119); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29121 = 12'h591 == _T_837 ? $signed(7'sh5) : $signed(_GEN_29120); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29122 = 12'h592 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29121); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29123 = 12'h593 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29122); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29124 = 12'h594 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29123); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29125 = 12'h595 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29124); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29126 = 12'h596 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29125); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29127 = 12'h597 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29126); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29128 = 12'h598 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29127); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29129 = 12'h599 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29128); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29130 = 12'h59a == _T_837 ? $signed(7'sh20) : $signed(_GEN_29129); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29131 = 12'h59b == _T_837 ? $signed(7'sh20) : $signed(_GEN_29130); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29132 = 12'h59c == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29131); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29133 = 12'h59d == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29132); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29134 = 12'h59e == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29133); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29135 = 12'h59f == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29134); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29136 = 12'h5a0 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29135); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29137 = 12'h5a1 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29136); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29138 = 12'h5a2 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29137); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29139 = 12'h5a3 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29138); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29140 = 12'h5a4 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29139); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29141 = 12'h5a5 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29140); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29142 = 12'h5a6 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29141); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29143 = 12'h5a7 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29142); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29144 = 12'h5a8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29143); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29145 = 12'h5a9 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29144); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29146 = 12'h5aa == _T_837 ? $signed(7'sh15) : $signed(_GEN_29145); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29147 = 12'h5ab == _T_837 ? $signed(7'sh14) : $signed(_GEN_29146); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29148 = 12'h5ac == _T_837 ? $signed(7'sh14) : $signed(_GEN_29147); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29149 = 12'h5ad == _T_837 ? $signed(7'sh13) : $signed(_GEN_29148); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29150 = 12'h5ae == _T_837 ? $signed(7'sh12) : $signed(_GEN_29149); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29151 = 12'h5af == _T_837 ? $signed(7'sh11) : $signed(_GEN_29150); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29152 = 12'h5b0 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29151); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29153 = 12'h5b1 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29152); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29154 = 12'h5b2 == _T_837 ? $signed(7'shf) : $signed(_GEN_29153); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29155 = 12'h5b3 == _T_837 ? $signed(7'shf) : $signed(_GEN_29154); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29156 = 12'h5b4 == _T_837 ? $signed(7'she) : $signed(_GEN_29155); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29157 = 12'h5b5 == _T_837 ? $signed(7'shd) : $signed(_GEN_29156); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29158 = 12'h5b6 == _T_837 ? $signed(7'shc) : $signed(_GEN_29157); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29159 = 12'h5b7 == _T_837 ? $signed(7'shc) : $signed(_GEN_29158); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29160 = 12'h5b8 == _T_837 ? $signed(7'shb) : $signed(_GEN_29159); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29161 = 12'h5b9 == _T_837 ? $signed(7'sha) : $signed(_GEN_29160); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29162 = 12'h5ba == _T_837 ? $signed(7'sha) : $signed(_GEN_29161); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29163 = 12'h5bb == _T_837 ? $signed(7'sh9) : $signed(_GEN_29162); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29164 = 12'h5bc == _T_837 ? $signed(7'sh8) : $signed(_GEN_29163); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29165 = 12'h5bd == _T_837 ? $signed(7'sh8) : $signed(_GEN_29164); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29166 = 12'h5be == _T_837 ? $signed(7'sh7) : $signed(_GEN_29165); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29167 = 12'h5bf == _T_837 ? $signed(7'sh6) : $signed(_GEN_29166); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29168 = 12'h5c0 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29167); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29169 = 12'h5c1 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29168); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29170 = 12'h5c2 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29169); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29171 = 12'h5c3 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29170); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29172 = 12'h5c4 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29171); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29173 = 12'h5c5 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29172); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29174 = 12'h5c6 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29173); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29175 = 12'h5c7 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29174); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29176 = 12'h5c8 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29175); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29177 = 12'h5c9 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29176); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29178 = 12'h5ca == _T_837 ? $signed(7'sh20) : $signed(_GEN_29177); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29179 = 12'h5cb == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29178); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29180 = 12'h5cc == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29179); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29181 = 12'h5cd == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29180); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29182 = 12'h5ce == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29181); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29183 = 12'h5cf == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29182); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29184 = 12'h5d0 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29183); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29185 = 12'h5d1 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29184); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29186 = 12'h5d2 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29185); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29187 = 12'h5d3 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29186); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29188 = 12'h5d4 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29187); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29189 = 12'h5d5 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29188); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29190 = 12'h5d6 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29189); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29191 = 12'h5d7 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29190); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29192 = 12'h5d8 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29191); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29193 = 12'h5d9 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29192); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29194 = 12'h5da == _T_837 ? $signed(7'sh14) : $signed(_GEN_29193); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29195 = 12'h5db == _T_837 ? $signed(7'sh14) : $signed(_GEN_29194); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29196 = 12'h5dc == _T_837 ? $signed(7'sh13) : $signed(_GEN_29195); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29197 = 12'h5dd == _T_837 ? $signed(7'sh12) : $signed(_GEN_29196); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29198 = 12'h5de == _T_837 ? $signed(7'sh11) : $signed(_GEN_29197); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29199 = 12'h5df == _T_837 ? $signed(7'sh11) : $signed(_GEN_29198); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29200 = 12'h5e0 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29199); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29201 = 12'h5e1 == _T_837 ? $signed(7'shf) : $signed(_GEN_29200); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29202 = 12'h5e2 == _T_837 ? $signed(7'shf) : $signed(_GEN_29201); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29203 = 12'h5e3 == _T_837 ? $signed(7'she) : $signed(_GEN_29202); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29204 = 12'h5e4 == _T_837 ? $signed(7'shd) : $signed(_GEN_29203); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29205 = 12'h5e5 == _T_837 ? $signed(7'shc) : $signed(_GEN_29204); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29206 = 12'h5e6 == _T_837 ? $signed(7'shc) : $signed(_GEN_29205); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29207 = 12'h5e7 == _T_837 ? $signed(7'shb) : $signed(_GEN_29206); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29208 = 12'h5e8 == _T_837 ? $signed(7'sha) : $signed(_GEN_29207); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29209 = 12'h5e9 == _T_837 ? $signed(7'sha) : $signed(_GEN_29208); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29210 = 12'h5ea == _T_837 ? $signed(7'sh9) : $signed(_GEN_29209); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29211 = 12'h5eb == _T_837 ? $signed(7'sh8) : $signed(_GEN_29210); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29212 = 12'h5ec == _T_837 ? $signed(7'sh8) : $signed(_GEN_29211); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29213 = 12'h5ed == _T_837 ? $signed(7'sh7) : $signed(_GEN_29212); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29214 = 12'h5ee == _T_837 ? $signed(7'sh27) : $signed(_GEN_29213); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29215 = 12'h5ef == _T_837 ? $signed(7'sh27) : $signed(_GEN_29214); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29216 = 12'h5f0 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29215); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29217 = 12'h5f1 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29216); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29218 = 12'h5f2 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29217); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29219 = 12'h5f3 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29218); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29220 = 12'h5f4 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29219); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29221 = 12'h5f5 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29220); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29222 = 12'h5f6 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29221); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29223 = 12'h5f7 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29222); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29224 = 12'h5f8 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29223); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29225 = 12'h5f9 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29224); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29226 = 12'h5fa == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29225); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29227 = 12'h5fb == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29226); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29228 = 12'h5fc == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29227); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29229 = 12'h5fd == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29228); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29230 = 12'h5fe == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29229); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29231 = 12'h5ff == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29230); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29232 = 12'h600 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29231); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29233 = 12'h601 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29232); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29234 = 12'h602 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29233); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29235 = 12'h603 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29234); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29236 = 12'h604 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29235); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29237 = 12'h605 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29236); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29238 = 12'h606 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29237); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29239 = 12'h607 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29238); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29240 = 12'h608 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29239); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29241 = 12'h609 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29240); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29242 = 12'h60a == _T_837 ? $signed(7'sh14) : $signed(_GEN_29241); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29243 = 12'h60b == _T_837 ? $signed(7'sh13) : $signed(_GEN_29242); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29244 = 12'h60c == _T_837 ? $signed(7'sh12) : $signed(_GEN_29243); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29245 = 12'h60d == _T_837 ? $signed(7'sh11) : $signed(_GEN_29244); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29246 = 12'h60e == _T_837 ? $signed(7'sh11) : $signed(_GEN_29245); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29247 = 12'h60f == _T_837 ? $signed(7'sh10) : $signed(_GEN_29246); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29248 = 12'h610 == _T_837 ? $signed(7'shf) : $signed(_GEN_29247); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29249 = 12'h611 == _T_837 ? $signed(7'shf) : $signed(_GEN_29248); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29250 = 12'h612 == _T_837 ? $signed(7'she) : $signed(_GEN_29249); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29251 = 12'h613 == _T_837 ? $signed(7'shd) : $signed(_GEN_29250); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29252 = 12'h614 == _T_837 ? $signed(7'shc) : $signed(_GEN_29251); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29253 = 12'h615 == _T_837 ? $signed(7'shc) : $signed(_GEN_29252); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29254 = 12'h616 == _T_837 ? $signed(7'shb) : $signed(_GEN_29253); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29255 = 12'h617 == _T_837 ? $signed(7'sha) : $signed(_GEN_29254); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29256 = 12'h618 == _T_837 ? $signed(7'sha) : $signed(_GEN_29255); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29257 = 12'h619 == _T_837 ? $signed(7'sh9) : $signed(_GEN_29256); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29258 = 12'h61a == _T_837 ? $signed(7'sh8) : $signed(_GEN_29257); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29259 = 12'h61b == _T_837 ? $signed(7'sh8) : $signed(_GEN_29258); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29260 = 12'h61c == _T_837 ? $signed(7'sh28) : $signed(_GEN_29259); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29261 = 12'h61d == _T_837 ? $signed(7'sh27) : $signed(_GEN_29260); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29262 = 12'h61e == _T_837 ? $signed(7'sh27) : $signed(_GEN_29261); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29263 = 12'h61f == _T_837 ? $signed(7'sh26) : $signed(_GEN_29262); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29264 = 12'h620 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29263); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29265 = 12'h621 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29264); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29266 = 12'h622 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29265); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29267 = 12'h623 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29266); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29268 = 12'h624 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29267); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29269 = 12'h625 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29268); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29270 = 12'h626 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29269); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29271 = 12'h627 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29270); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29272 = 12'h628 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29271); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29273 = 12'h629 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29272); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29274 = 12'h62a == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29273); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29275 = 12'h62b == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29274); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29276 = 12'h62c == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29275); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29277 = 12'h62d == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29276); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29278 = 12'h62e == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29277); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29279 = 12'h62f == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29278); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29280 = 12'h630 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29279); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29281 = 12'h631 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29280); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29282 = 12'h632 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29281); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29283 = 12'h633 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29282); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29284 = 12'h634 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29283); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29285 = 12'h635 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29284); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29286 = 12'h636 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29285); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29287 = 12'h637 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29286); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29288 = 12'h638 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29287); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29289 = 12'h639 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29288); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29290 = 12'h63a == _T_837 ? $signed(7'sh13) : $signed(_GEN_29289); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29291 = 12'h63b == _T_837 ? $signed(7'sh12) : $signed(_GEN_29290); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29292 = 12'h63c == _T_837 ? $signed(7'sh11) : $signed(_GEN_29291); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29293 = 12'h63d == _T_837 ? $signed(7'sh11) : $signed(_GEN_29292); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29294 = 12'h63e == _T_837 ? $signed(7'sh10) : $signed(_GEN_29293); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29295 = 12'h63f == _T_837 ? $signed(7'shf) : $signed(_GEN_29294); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29296 = 12'h640 == _T_837 ? $signed(7'shf) : $signed(_GEN_29295); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29297 = 12'h641 == _T_837 ? $signed(7'she) : $signed(_GEN_29296); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29298 = 12'h642 == _T_837 ? $signed(7'shd) : $signed(_GEN_29297); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29299 = 12'h643 == _T_837 ? $signed(7'shc) : $signed(_GEN_29298); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29300 = 12'h644 == _T_837 ? $signed(7'shc) : $signed(_GEN_29299); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29301 = 12'h645 == _T_837 ? $signed(7'shb) : $signed(_GEN_29300); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29302 = 12'h646 == _T_837 ? $signed(7'sha) : $signed(_GEN_29301); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29303 = 12'h647 == _T_837 ? $signed(7'sha) : $signed(_GEN_29302); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29304 = 12'h648 == _T_837 ? $signed(7'sh9) : $signed(_GEN_29303); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29305 = 12'h649 == _T_837 ? $signed(7'sh8) : $signed(_GEN_29304); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29306 = 12'h64a == _T_837 ? $signed(7'sh29) : $signed(_GEN_29305); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29307 = 12'h64b == _T_837 ? $signed(7'sh28) : $signed(_GEN_29306); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29308 = 12'h64c == _T_837 ? $signed(7'sh27) : $signed(_GEN_29307); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29309 = 12'h64d == _T_837 ? $signed(7'sh27) : $signed(_GEN_29308); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29310 = 12'h64e == _T_837 ? $signed(7'sh26) : $signed(_GEN_29309); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29311 = 12'h64f == _T_837 ? $signed(7'sh25) : $signed(_GEN_29310); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29312 = 12'h650 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29311); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29313 = 12'h651 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29312); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29314 = 12'h652 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29313); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29315 = 12'h653 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29314); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29316 = 12'h654 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29315); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29317 = 12'h655 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29316); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29318 = 12'h656 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29317); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29319 = 12'h657 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29318); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29320 = 12'h658 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29319); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29321 = 12'h659 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29320); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29322 = 12'h65a == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29321); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29323 = 12'h65b == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29322); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29324 = 12'h65c == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29323); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29325 = 12'h65d == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29324); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29326 = 12'h65e == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29325); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29327 = 12'h65f == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29326); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29328 = 12'h660 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29327); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29329 = 12'h661 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29328); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29330 = 12'h662 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29329); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29331 = 12'h663 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29330); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29332 = 12'h664 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29331); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29333 = 12'h665 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29332); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29334 = 12'h666 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29333); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29335 = 12'h667 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29334); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29336 = 12'h668 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29335); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29337 = 12'h669 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29336); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29338 = 12'h66a == _T_837 ? $signed(7'sh12) : $signed(_GEN_29337); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29339 = 12'h66b == _T_837 ? $signed(7'sh11) : $signed(_GEN_29338); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29340 = 12'h66c == _T_837 ? $signed(7'sh11) : $signed(_GEN_29339); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29341 = 12'h66d == _T_837 ? $signed(7'sh10) : $signed(_GEN_29340); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29342 = 12'h66e == _T_837 ? $signed(7'shf) : $signed(_GEN_29341); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29343 = 12'h66f == _T_837 ? $signed(7'shf) : $signed(_GEN_29342); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29344 = 12'h670 == _T_837 ? $signed(7'she) : $signed(_GEN_29343); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29345 = 12'h671 == _T_837 ? $signed(7'shd) : $signed(_GEN_29344); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29346 = 12'h672 == _T_837 ? $signed(7'shc) : $signed(_GEN_29345); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29347 = 12'h673 == _T_837 ? $signed(7'shc) : $signed(_GEN_29346); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29348 = 12'h674 == _T_837 ? $signed(7'shb) : $signed(_GEN_29347); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29349 = 12'h675 == _T_837 ? $signed(7'sha) : $signed(_GEN_29348); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29350 = 12'h676 == _T_837 ? $signed(7'sha) : $signed(_GEN_29349); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29351 = 12'h677 == _T_837 ? $signed(7'sh9) : $signed(_GEN_29350); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29352 = 12'h678 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29351); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29353 = 12'h679 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29352); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29354 = 12'h67a == _T_837 ? $signed(7'sh28) : $signed(_GEN_29353); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29355 = 12'h67b == _T_837 ? $signed(7'sh27) : $signed(_GEN_29354); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29356 = 12'h67c == _T_837 ? $signed(7'sh27) : $signed(_GEN_29355); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29357 = 12'h67d == _T_837 ? $signed(7'sh26) : $signed(_GEN_29356); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29358 = 12'h67e == _T_837 ? $signed(7'sh25) : $signed(_GEN_29357); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29359 = 12'h67f == _T_837 ? $signed(7'sh25) : $signed(_GEN_29358); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29360 = 12'h680 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29359); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29361 = 12'h681 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29360); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29362 = 12'h682 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29361); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29363 = 12'h683 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29362); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29364 = 12'h684 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29363); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29365 = 12'h685 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29364); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29366 = 12'h686 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29365); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29367 = 12'h687 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29366); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29368 = 12'h688 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29367); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29369 = 12'h689 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29368); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29370 = 12'h68a == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29369); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29371 = 12'h68b == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29370); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29372 = 12'h68c == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29371); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29373 = 12'h68d == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29372); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29374 = 12'h68e == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29373); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29375 = 12'h68f == _T_837 ? $signed(7'sh19) : $signed(_GEN_29374); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29376 = 12'h690 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29375); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29377 = 12'h691 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29376); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29378 = 12'h692 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29377); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29379 = 12'h693 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29378); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29380 = 12'h694 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29379); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29381 = 12'h695 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29380); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29382 = 12'h696 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29381); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29383 = 12'h697 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29382); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29384 = 12'h698 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29383); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29385 = 12'h699 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29384); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29386 = 12'h69a == _T_837 ? $signed(7'sh11) : $signed(_GEN_29385); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29387 = 12'h69b == _T_837 ? $signed(7'sh11) : $signed(_GEN_29386); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29388 = 12'h69c == _T_837 ? $signed(7'sh10) : $signed(_GEN_29387); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29389 = 12'h69d == _T_837 ? $signed(7'shf) : $signed(_GEN_29388); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29390 = 12'h69e == _T_837 ? $signed(7'shf) : $signed(_GEN_29389); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29391 = 12'h69f == _T_837 ? $signed(7'she) : $signed(_GEN_29390); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29392 = 12'h6a0 == _T_837 ? $signed(7'shd) : $signed(_GEN_29391); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29393 = 12'h6a1 == _T_837 ? $signed(7'shc) : $signed(_GEN_29392); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29394 = 12'h6a2 == _T_837 ? $signed(7'shc) : $signed(_GEN_29393); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29395 = 12'h6a3 == _T_837 ? $signed(7'shb) : $signed(_GEN_29394); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29396 = 12'h6a4 == _T_837 ? $signed(7'sha) : $signed(_GEN_29395); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29397 = 12'h6a5 == _T_837 ? $signed(7'sha) : $signed(_GEN_29396); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29398 = 12'h6a6 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29397); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29399 = 12'h6a7 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29398); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29400 = 12'h6a8 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29399); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29401 = 12'h6a9 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29400); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29402 = 12'h6aa == _T_837 ? $signed(7'sh27) : $signed(_GEN_29401); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29403 = 12'h6ab == _T_837 ? $signed(7'sh27) : $signed(_GEN_29402); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29404 = 12'h6ac == _T_837 ? $signed(7'sh26) : $signed(_GEN_29403); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29405 = 12'h6ad == _T_837 ? $signed(7'sh25) : $signed(_GEN_29404); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29406 = 12'h6ae == _T_837 ? $signed(7'sh25) : $signed(_GEN_29405); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29407 = 12'h6af == _T_837 ? $signed(7'sh24) : $signed(_GEN_29406); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29408 = 12'h6b0 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29407); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29409 = 12'h6b1 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29408); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29410 = 12'h6b2 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29409); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29411 = 12'h6b3 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29410); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29412 = 12'h6b4 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29411); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29413 = 12'h6b5 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29412); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29414 = 12'h6b6 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29413); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29415 = 12'h6b7 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29414); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29416 = 12'h6b8 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29415); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29417 = 12'h6b9 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29416); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29418 = 12'h6ba == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29417); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29419 = 12'h6bb == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29418); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29420 = 12'h6bc == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29419); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29421 = 12'h6bd == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29420); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29422 = 12'h6be == _T_837 ? $signed(7'sh19) : $signed(_GEN_29421); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29423 = 12'h6bf == _T_837 ? $signed(7'sh18) : $signed(_GEN_29422); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29424 = 12'h6c0 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29423); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29425 = 12'h6c1 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29424); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29426 = 12'h6c2 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29425); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29427 = 12'h6c3 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29426); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29428 = 12'h6c4 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29427); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29429 = 12'h6c5 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29428); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29430 = 12'h6c6 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29429); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29431 = 12'h6c7 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29430); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29432 = 12'h6c8 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29431); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29433 = 12'h6c9 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29432); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29434 = 12'h6ca == _T_837 ? $signed(7'sh11) : $signed(_GEN_29433); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29435 = 12'h6cb == _T_837 ? $signed(7'sh10) : $signed(_GEN_29434); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29436 = 12'h6cc == _T_837 ? $signed(7'shf) : $signed(_GEN_29435); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29437 = 12'h6cd == _T_837 ? $signed(7'shf) : $signed(_GEN_29436); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29438 = 12'h6ce == _T_837 ? $signed(7'she) : $signed(_GEN_29437); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29439 = 12'h6cf == _T_837 ? $signed(7'shd) : $signed(_GEN_29438); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29440 = 12'h6d0 == _T_837 ? $signed(7'shc) : $signed(_GEN_29439); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29441 = 12'h6d1 == _T_837 ? $signed(7'shc) : $signed(_GEN_29440); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29442 = 12'h6d2 == _T_837 ? $signed(7'shb) : $signed(_GEN_29441); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29443 = 12'h6d3 == _T_837 ? $signed(7'sha) : $signed(_GEN_29442); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29444 = 12'h6d4 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29443); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29445 = 12'h6d5 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29444); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29446 = 12'h6d6 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29445); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29447 = 12'h6d7 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29446); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29448 = 12'h6d8 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29447); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29449 = 12'h6d9 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29448); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29450 = 12'h6da == _T_837 ? $signed(7'sh27) : $signed(_GEN_29449); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29451 = 12'h6db == _T_837 ? $signed(7'sh26) : $signed(_GEN_29450); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29452 = 12'h6dc == _T_837 ? $signed(7'sh25) : $signed(_GEN_29451); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29453 = 12'h6dd == _T_837 ? $signed(7'sh25) : $signed(_GEN_29452); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29454 = 12'h6de == _T_837 ? $signed(7'sh24) : $signed(_GEN_29453); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29455 = 12'h6df == _T_837 ? $signed(7'sh23) : $signed(_GEN_29454); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29456 = 12'h6e0 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29455); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29457 = 12'h6e1 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29456); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29458 = 12'h6e2 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29457); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29459 = 12'h6e3 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29458); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29460 = 12'h6e4 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29459); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29461 = 12'h6e5 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29460); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29462 = 12'h6e6 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29461); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29463 = 12'h6e7 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29462); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29464 = 12'h6e8 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29463); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29465 = 12'h6e9 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29464); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29466 = 12'h6ea == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29465); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29467 = 12'h6eb == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29466); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29468 = 12'h6ec == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29467); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29469 = 12'h6ed == _T_837 ? $signed(7'sh19) : $signed(_GEN_29468); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29470 = 12'h6ee == _T_837 ? $signed(7'sh18) : $signed(_GEN_29469); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29471 = 12'h6ef == _T_837 ? $signed(7'sh18) : $signed(_GEN_29470); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29472 = 12'h6f0 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29471); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29473 = 12'h6f1 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29472); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29474 = 12'h6f2 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29473); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29475 = 12'h6f3 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29474); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29476 = 12'h6f4 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29475); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29477 = 12'h6f5 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29476); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29478 = 12'h6f6 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29477); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29479 = 12'h6f7 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29478); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29480 = 12'h6f8 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29479); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29481 = 12'h6f9 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29480); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29482 = 12'h6fa == _T_837 ? $signed(7'sh10) : $signed(_GEN_29481); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29483 = 12'h6fb == _T_837 ? $signed(7'shf) : $signed(_GEN_29482); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29484 = 12'h6fc == _T_837 ? $signed(7'shf) : $signed(_GEN_29483); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29485 = 12'h6fd == _T_837 ? $signed(7'she) : $signed(_GEN_29484); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29486 = 12'h6fe == _T_837 ? $signed(7'shd) : $signed(_GEN_29485); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29487 = 12'h6ff == _T_837 ? $signed(7'shc) : $signed(_GEN_29486); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29488 = 12'h700 == _T_837 ? $signed(7'shc) : $signed(_GEN_29487); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29489 = 12'h701 == _T_837 ? $signed(7'shb) : $signed(_GEN_29488); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29490 = 12'h702 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29489); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29491 = 12'h703 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29490); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29492 = 12'h704 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29491); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29493 = 12'h705 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29492); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29494 = 12'h706 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29493); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29495 = 12'h707 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29494); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29496 = 12'h708 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29495); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29497 = 12'h709 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29496); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29498 = 12'h70a == _T_837 ? $signed(7'sh26) : $signed(_GEN_29497); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29499 = 12'h70b == _T_837 ? $signed(7'sh25) : $signed(_GEN_29498); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29500 = 12'h70c == _T_837 ? $signed(7'sh25) : $signed(_GEN_29499); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29501 = 12'h70d == _T_837 ? $signed(7'sh24) : $signed(_GEN_29500); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29502 = 12'h70e == _T_837 ? $signed(7'sh23) : $signed(_GEN_29501); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29503 = 12'h70f == _T_837 ? $signed(7'sh22) : $signed(_GEN_29502); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29504 = 12'h710 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29503); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29505 = 12'h711 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29504); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29506 = 12'h712 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29505); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29507 = 12'h713 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29506); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29508 = 12'h714 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29507); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29509 = 12'h715 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29508); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29510 = 12'h716 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29509); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29511 = 12'h717 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29510); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29512 = 12'h718 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29511); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29513 = 12'h719 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29512); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29514 = 12'h71a == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29513); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29515 = 12'h71b == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29514); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29516 = 12'h71c == _T_837 ? $signed(7'sh19) : $signed(_GEN_29515); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29517 = 12'h71d == _T_837 ? $signed(7'sh18) : $signed(_GEN_29516); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29518 = 12'h71e == _T_837 ? $signed(7'sh18) : $signed(_GEN_29517); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29519 = 12'h71f == _T_837 ? $signed(7'sh17) : $signed(_GEN_29518); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29520 = 12'h720 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29519); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29521 = 12'h721 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29520); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29522 = 12'h722 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29521); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29523 = 12'h723 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29522); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29524 = 12'h724 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29523); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29525 = 12'h725 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29524); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29526 = 12'h726 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29525); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29527 = 12'h727 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29526); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29528 = 12'h728 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29527); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29529 = 12'h729 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29528); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29530 = 12'h72a == _T_837 ? $signed(7'shf) : $signed(_GEN_29529); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29531 = 12'h72b == _T_837 ? $signed(7'shf) : $signed(_GEN_29530); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29532 = 12'h72c == _T_837 ? $signed(7'she) : $signed(_GEN_29531); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29533 = 12'h72d == _T_837 ? $signed(7'shd) : $signed(_GEN_29532); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29534 = 12'h72e == _T_837 ? $signed(7'shc) : $signed(_GEN_29533); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29535 = 12'h72f == _T_837 ? $signed(7'shc) : $signed(_GEN_29534); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29536 = 12'h730 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29535); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29537 = 12'h731 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29536); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29538 = 12'h732 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29537); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29539 = 12'h733 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29538); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29540 = 12'h734 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29539); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29541 = 12'h735 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29540); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29542 = 12'h736 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29541); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29543 = 12'h737 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29542); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29544 = 12'h738 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29543); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29545 = 12'h739 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29544); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29546 = 12'h73a == _T_837 ? $signed(7'sh25) : $signed(_GEN_29545); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29547 = 12'h73b == _T_837 ? $signed(7'sh25) : $signed(_GEN_29546); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29548 = 12'h73c == _T_837 ? $signed(7'sh24) : $signed(_GEN_29547); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29549 = 12'h73d == _T_837 ? $signed(7'sh23) : $signed(_GEN_29548); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29550 = 12'h73e == _T_837 ? $signed(7'sh22) : $signed(_GEN_29549); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29551 = 12'h73f == _T_837 ? $signed(7'sh22) : $signed(_GEN_29550); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29552 = 12'h740 == _T_837 ? $signed(7'sh21) : $signed(_GEN_29551); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29553 = 12'h741 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29552); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29554 = 12'h742 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29553); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29555 = 12'h743 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29554); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29556 = 12'h744 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29555); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29557 = 12'h745 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29556); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29558 = 12'h746 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29557); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29559 = 12'h747 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29558); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29560 = 12'h748 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29559); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29561 = 12'h749 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29560); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29562 = 12'h74a == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29561); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29563 = 12'h74b == _T_837 ? $signed(7'sh19) : $signed(_GEN_29562); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29564 = 12'h74c == _T_837 ? $signed(7'sh18) : $signed(_GEN_29563); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29565 = 12'h74d == _T_837 ? $signed(7'sh18) : $signed(_GEN_29564); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29566 = 12'h74e == _T_837 ? $signed(7'sh17) : $signed(_GEN_29565); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29567 = 12'h74f == _T_837 ? $signed(7'sh16) : $signed(_GEN_29566); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29568 = 12'h750 == _T_837 ? $signed(7'sh16) : $signed(_GEN_29567); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29569 = 12'h751 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29568); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29570 = 12'h752 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29569); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29571 = 12'h753 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29570); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29572 = 12'h754 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29571); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29573 = 12'h755 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29572); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29574 = 12'h756 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29573); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29575 = 12'h757 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29574); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29576 = 12'h758 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29575); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29577 = 12'h759 == _T_837 ? $signed(7'shf) : $signed(_GEN_29576); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29578 = 12'h75a == _T_837 ? $signed(7'shf) : $signed(_GEN_29577); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29579 = 12'h75b == _T_837 ? $signed(7'she) : $signed(_GEN_29578); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29580 = 12'h75c == _T_837 ? $signed(7'shd) : $signed(_GEN_29579); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29581 = 12'h75d == _T_837 ? $signed(7'shc) : $signed(_GEN_29580); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29582 = 12'h75e == _T_837 ? $signed(7'sh2d) : $signed(_GEN_29581); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29583 = 12'h75f == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29582); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29584 = 12'h760 == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29583); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29585 = 12'h761 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29584); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29586 = 12'h762 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29585); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29587 = 12'h763 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29586); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29588 = 12'h764 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29587); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29589 = 12'h765 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29588); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29590 = 12'h766 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29589); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29591 = 12'h767 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29590); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29592 = 12'h768 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29591); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29593 = 12'h769 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29592); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29594 = 12'h76a == _T_837 ? $signed(7'sh25) : $signed(_GEN_29593); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29595 = 12'h76b == _T_837 ? $signed(7'sh24) : $signed(_GEN_29594); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29596 = 12'h76c == _T_837 ? $signed(7'sh23) : $signed(_GEN_29595); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29597 = 12'h76d == _T_837 ? $signed(7'sh22) : $signed(_GEN_29596); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29598 = 12'h76e == _T_837 ? $signed(7'sh22) : $signed(_GEN_29597); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29599 = 12'h76f == _T_837 ? $signed(7'sh21) : $signed(_GEN_29598); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29600 = 12'h770 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29599); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29601 = 12'h771 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29600); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29602 = 12'h772 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29601); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29603 = 12'h773 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29602); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29604 = 12'h774 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29603); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29605 = 12'h775 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29604); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29606 = 12'h776 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29605); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29607 = 12'h777 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29606); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29608 = 12'h778 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29607); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29609 = 12'h779 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29608); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29610 = 12'h77a == _T_837 ? $signed(7'sh19) : $signed(_GEN_29609); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29611 = 12'h77b == _T_837 ? $signed(7'sh18) : $signed(_GEN_29610); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29612 = 12'h77c == _T_837 ? $signed(7'sh18) : $signed(_GEN_29611); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29613 = 12'h77d == _T_837 ? $signed(7'sh17) : $signed(_GEN_29612); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29614 = 12'h77e == _T_837 ? $signed(7'sh16) : $signed(_GEN_29613); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29615 = 12'h77f == _T_837 ? $signed(7'sh16) : $signed(_GEN_29614); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29616 = 12'h780 == _T_837 ? $signed(7'sh15) : $signed(_GEN_29615); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29617 = 12'h781 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29616); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29618 = 12'h782 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29617); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29619 = 12'h783 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29618); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29620 = 12'h784 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29619); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29621 = 12'h785 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29620); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29622 = 12'h786 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29621); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29623 = 12'h787 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29622); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29624 = 12'h788 == _T_837 ? $signed(7'shf) : $signed(_GEN_29623); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29625 = 12'h789 == _T_837 ? $signed(7'shf) : $signed(_GEN_29624); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29626 = 12'h78a == _T_837 ? $signed(7'she) : $signed(_GEN_29625); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29627 = 12'h78b == _T_837 ? $signed(7'shd) : $signed(_GEN_29626); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29628 = 12'h78c == _T_837 ? $signed(7'sh2e) : $signed(_GEN_29627); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29629 = 12'h78d == _T_837 ? $signed(7'sh2d) : $signed(_GEN_29628); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29630 = 12'h78e == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29629); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29631 = 12'h78f == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29630); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29632 = 12'h790 == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29631); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29633 = 12'h791 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29632); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29634 = 12'h792 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29633); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29635 = 12'h793 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29634); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29636 = 12'h794 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29635); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29637 = 12'h795 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29636); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29638 = 12'h796 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29637); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29639 = 12'h797 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29638); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29640 = 12'h798 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29639); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29641 = 12'h799 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29640); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29642 = 12'h79a == _T_837 ? $signed(7'sh24) : $signed(_GEN_29641); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29643 = 12'h79b == _T_837 ? $signed(7'sh23) : $signed(_GEN_29642); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29644 = 12'h79c == _T_837 ? $signed(7'sh22) : $signed(_GEN_29643); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29645 = 12'h79d == _T_837 ? $signed(7'sh22) : $signed(_GEN_29644); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29646 = 12'h79e == _T_837 ? $signed(7'sh21) : $signed(_GEN_29645); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29647 = 12'h79f == _T_837 ? $signed(7'sh20) : $signed(_GEN_29646); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29648 = 12'h7a0 == _T_837 ? $signed(7'sh20) : $signed(_GEN_29647); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29649 = 12'h7a1 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29648); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29650 = 12'h7a2 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29649); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29651 = 12'h7a3 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29650); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29652 = 12'h7a4 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29651); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29653 = 12'h7a5 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29652); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29654 = 12'h7a6 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29653); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29655 = 12'h7a7 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29654); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29656 = 12'h7a8 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29655); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29657 = 12'h7a9 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29656); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29658 = 12'h7aa == _T_837 ? $signed(7'sh18) : $signed(_GEN_29657); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29659 = 12'h7ab == _T_837 ? $signed(7'sh18) : $signed(_GEN_29658); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29660 = 12'h7ac == _T_837 ? $signed(7'sh17) : $signed(_GEN_29659); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29661 = 12'h7ad == _T_837 ? $signed(7'sh16) : $signed(_GEN_29660); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29662 = 12'h7ae == _T_837 ? $signed(7'sh16) : $signed(_GEN_29661); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29663 = 12'h7af == _T_837 ? $signed(7'sh15) : $signed(_GEN_29662); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29664 = 12'h7b0 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29663); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29665 = 12'h7b1 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29664); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29666 = 12'h7b2 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29665); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29667 = 12'h7b3 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29666); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29668 = 12'h7b4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29667); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29669 = 12'h7b5 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29668); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29670 = 12'h7b6 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29669); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29671 = 12'h7b7 == _T_837 ? $signed(7'shf) : $signed(_GEN_29670); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29672 = 12'h7b8 == _T_837 ? $signed(7'shf) : $signed(_GEN_29671); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29673 = 12'h7b9 == _T_837 ? $signed(7'she) : $signed(_GEN_29672); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29674 = 12'h7ba == _T_837 ? $signed(7'sh2e) : $signed(_GEN_29673); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29675 = 12'h7bb == _T_837 ? $signed(7'sh2e) : $signed(_GEN_29674); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29676 = 12'h7bc == _T_837 ? $signed(7'sh2d) : $signed(_GEN_29675); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29677 = 12'h7bd == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29676); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29678 = 12'h7be == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29677); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29679 = 12'h7bf == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29678); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29680 = 12'h7c0 == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29679); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29681 = 12'h7c1 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29680); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29682 = 12'h7c2 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29681); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29683 = 12'h7c3 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29682); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29684 = 12'h7c4 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29683); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29685 = 12'h7c5 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29684); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29686 = 12'h7c6 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29685); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29687 = 12'h7c7 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29686); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29688 = 12'h7c8 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29687); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29689 = 12'h7c9 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29688); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29690 = 12'h7ca == _T_837 ? $signed(7'sh23) : $signed(_GEN_29689); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29691 = 12'h7cb == _T_837 ? $signed(7'sh22) : $signed(_GEN_29690); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29692 = 12'h7cc == _T_837 ? $signed(7'sh22) : $signed(_GEN_29691); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29693 = 12'h7cd == _T_837 ? $signed(7'sh21) : $signed(_GEN_29692); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29694 = 12'h7ce == _T_837 ? $signed(7'sh20) : $signed(_GEN_29693); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29695 = 12'h7cf == _T_837 ? $signed(7'sh20) : $signed(_GEN_29694); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29696 = 12'h7d0 == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29695); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29697 = 12'h7d1 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29696); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29698 = 12'h7d2 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29697); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29699 = 12'h7d3 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29698); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29700 = 12'h7d4 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29699); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29701 = 12'h7d5 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29700); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29702 = 12'h7d6 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29701); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29703 = 12'h7d7 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29702); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29704 = 12'h7d8 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29703); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29705 = 12'h7d9 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29704); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29706 = 12'h7da == _T_837 ? $signed(7'sh18) : $signed(_GEN_29705); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29707 = 12'h7db == _T_837 ? $signed(7'sh17) : $signed(_GEN_29706); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29708 = 12'h7dc == _T_837 ? $signed(7'sh16) : $signed(_GEN_29707); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29709 = 12'h7dd == _T_837 ? $signed(7'sh16) : $signed(_GEN_29708); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29710 = 12'h7de == _T_837 ? $signed(7'sh15) : $signed(_GEN_29709); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29711 = 12'h7df == _T_837 ? $signed(7'sh14) : $signed(_GEN_29710); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29712 = 12'h7e0 == _T_837 ? $signed(7'sh14) : $signed(_GEN_29711); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29713 = 12'h7e1 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29712); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29714 = 12'h7e2 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29713); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29715 = 12'h7e3 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29714); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29716 = 12'h7e4 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29715); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29717 = 12'h7e5 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29716); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29718 = 12'h7e6 == _T_837 ? $signed(7'shf) : $signed(_GEN_29717); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29719 = 12'h7e7 == _T_837 ? $signed(7'shf) : $signed(_GEN_29718); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29720 = 12'h7e8 == _T_837 ? $signed(7'sh2f) : $signed(_GEN_29719); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29721 = 12'h7e9 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_29720); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29722 = 12'h7ea == _T_837 ? $signed(7'sh2e) : $signed(_GEN_29721); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29723 = 12'h7eb == _T_837 ? $signed(7'sh2d) : $signed(_GEN_29722); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29724 = 12'h7ec == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29723); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29725 = 12'h7ed == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29724); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29726 = 12'h7ee == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29725); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29727 = 12'h7ef == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29726); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29728 = 12'h7f0 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29727); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29729 = 12'h7f1 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29728); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29730 = 12'h7f2 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29729); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29731 = 12'h7f3 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29730); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29732 = 12'h7f4 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29731); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29733 = 12'h7f5 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29732); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29734 = 12'h7f6 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29733); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29735 = 12'h7f7 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29734); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29736 = 12'h7f8 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29735); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29737 = 12'h7f9 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29736); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29738 = 12'h7fa == _T_837 ? $signed(7'sh22) : $signed(_GEN_29737); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29739 = 12'h7fb == _T_837 ? $signed(7'sh22) : $signed(_GEN_29738); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29740 = 12'h7fc == _T_837 ? $signed(7'sh21) : $signed(_GEN_29739); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29741 = 12'h7fd == _T_837 ? $signed(7'sh20) : $signed(_GEN_29740); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29742 = 12'h7fe == _T_837 ? $signed(7'sh20) : $signed(_GEN_29741); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29743 = 12'h7ff == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29742); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29744 = 12'h800 == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29743); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29745 = 12'h801 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29744); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29746 = 12'h802 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29745); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29747 = 12'h803 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29746); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29748 = 12'h804 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29747); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29749 = 12'h805 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29748); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29750 = 12'h806 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29749); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29751 = 12'h807 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29750); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29752 = 12'h808 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29751); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29753 = 12'h809 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29752); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29754 = 12'h80a == _T_837 ? $signed(7'sh17) : $signed(_GEN_29753); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29755 = 12'h80b == _T_837 ? $signed(7'sh16) : $signed(_GEN_29754); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29756 = 12'h80c == _T_837 ? $signed(7'sh16) : $signed(_GEN_29755); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29757 = 12'h80d == _T_837 ? $signed(7'sh15) : $signed(_GEN_29756); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29758 = 12'h80e == _T_837 ? $signed(7'sh14) : $signed(_GEN_29757); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29759 = 12'h80f == _T_837 ? $signed(7'sh14) : $signed(_GEN_29758); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29760 = 12'h810 == _T_837 ? $signed(7'sh13) : $signed(_GEN_29759); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29761 = 12'h811 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29760); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29762 = 12'h812 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29761); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29763 = 12'h813 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29762); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29764 = 12'h814 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29763); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29765 = 12'h815 == _T_837 ? $signed(7'shf) : $signed(_GEN_29764); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29766 = 12'h816 == _T_837 ? $signed(7'sh30) : $signed(_GEN_29765); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29767 = 12'h817 == _T_837 ? $signed(7'sh2f) : $signed(_GEN_29766); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29768 = 12'h818 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_29767); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29769 = 12'h819 == _T_837 ? $signed(7'sh2e) : $signed(_GEN_29768); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29770 = 12'h81a == _T_837 ? $signed(7'sh2d) : $signed(_GEN_29769); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29771 = 12'h81b == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29770); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29772 = 12'h81c == _T_837 ? $signed(7'sh2c) : $signed(_GEN_29771); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29773 = 12'h81d == _T_837 ? $signed(7'sh2b) : $signed(_GEN_29772); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29774 = 12'h81e == _T_837 ? $signed(7'sh2a) : $signed(_GEN_29773); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29775 = 12'h81f == _T_837 ? $signed(7'sh29) : $signed(_GEN_29774); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29776 = 12'h820 == _T_837 ? $signed(7'sh29) : $signed(_GEN_29775); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29777 = 12'h821 == _T_837 ? $signed(7'sh28) : $signed(_GEN_29776); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29778 = 12'h822 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29777); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29779 = 12'h823 == _T_837 ? $signed(7'sh27) : $signed(_GEN_29778); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29780 = 12'h824 == _T_837 ? $signed(7'sh26) : $signed(_GEN_29779); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29781 = 12'h825 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29780); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29782 = 12'h826 == _T_837 ? $signed(7'sh25) : $signed(_GEN_29781); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29783 = 12'h827 == _T_837 ? $signed(7'sh24) : $signed(_GEN_29782); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29784 = 12'h828 == _T_837 ? $signed(7'sh23) : $signed(_GEN_29783); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29785 = 12'h829 == _T_837 ? $signed(7'sh22) : $signed(_GEN_29784); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29786 = 12'h82a == _T_837 ? $signed(7'sh22) : $signed(_GEN_29785); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29787 = 12'h82b == _T_837 ? $signed(7'sh21) : $signed(_GEN_29786); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29788 = 12'h82c == _T_837 ? $signed(7'sh20) : $signed(_GEN_29787); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29789 = 12'h82d == _T_837 ? $signed(7'sh20) : $signed(_GEN_29788); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29790 = 12'h82e == _T_837 ? $signed(7'sh1f) : $signed(_GEN_29789); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29791 = 12'h82f == _T_837 ? $signed(7'sh1e) : $signed(_GEN_29790); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29792 = 12'h830 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29791); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29793 = 12'h831 == _T_837 ? $signed(7'sh1d) : $signed(_GEN_29792); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29794 = 12'h832 == _T_837 ? $signed(7'sh1c) : $signed(_GEN_29793); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29795 = 12'h833 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29794); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29796 = 12'h834 == _T_837 ? $signed(7'sh1b) : $signed(_GEN_29795); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29797 = 12'h835 == _T_837 ? $signed(7'sh1a) : $signed(_GEN_29796); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29798 = 12'h836 == _T_837 ? $signed(7'sh19) : $signed(_GEN_29797); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29799 = 12'h837 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29798); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29800 = 12'h838 == _T_837 ? $signed(7'sh18) : $signed(_GEN_29799); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29801 = 12'h839 == _T_837 ? $signed(7'sh17) : $signed(_GEN_29800); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29802 = 12'h83a == _T_837 ? $signed(7'sh16) : $signed(_GEN_29801); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29803 = 12'h83b == _T_837 ? $signed(7'sh16) : $signed(_GEN_29802); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29804 = 12'h83c == _T_837 ? $signed(7'sh15) : $signed(_GEN_29803); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29805 = 12'h83d == _T_837 ? $signed(7'sh14) : $signed(_GEN_29804); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29806 = 12'h83e == _T_837 ? $signed(7'sh14) : $signed(_GEN_29805); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29807 = 12'h83f == _T_837 ? $signed(7'sh13) : $signed(_GEN_29806); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29808 = 12'h840 == _T_837 ? $signed(7'sh12) : $signed(_GEN_29807); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29809 = 12'h841 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29808); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29810 = 12'h842 == _T_837 ? $signed(7'sh11) : $signed(_GEN_29809); // @[GraphicEngineVGA.scala 322:24]
  wire [6:0] _GEN_29811 = 12'h843 == _T_837 ? $signed(7'sh10) : $signed(_GEN_29810); // @[GraphicEngineVGA.scala 322:24]
  wire [11:0] _T_839 = spriteRotationReg_6 ? $signed({{5{_GEN_29811[6]}},_GEN_29811}) : $signed(_T_832); // @[GraphicEngineVGA.scala 322:24]
  wire [10:0] inSpriteY_6 = _T_839[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire  _T_866 = $signed(_T_822) >= 12'sh0; // @[GraphicEngineVGA.scala 343:27]
  wire  _T_867 = $signed(_T_822) < 12'sh2e; // @[GraphicEngineVGA.scala 343:47]
  wire  _T_868 = _T_866 & _T_867; // @[GraphicEngineVGA.scala 343:35]
  wire  _T_869 = $signed(_T_832) >= 12'sh0; // @[GraphicEngineVGA.scala 344:27]
  wire  _T_870 = $signed(_T_832) < 12'sh2e; // @[GraphicEngineVGA.scala 344:47]
  wire  _T_871 = _T_869 & _T_870; // @[GraphicEngineVGA.scala 344:35]
  wire  _T_872 = _T_868 & _T_871; // @[GraphicEngineVGA.scala 345:32]
  wire  _T_873 = $signed(inSpriteX_6) >= 12'sh0; // @[GraphicEngineVGA.scala 347:31]
  wire  _T_874 = $signed(inSpriteX_6) < 12'sh20; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_875 = _T_873 & _T_874; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_876 = $signed(inSpriteY_6) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire  _T_877 = $signed(inSpriteY_6) < 11'sh20; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_878 = _T_876 & _T_877; // @[GraphicEngineVGA.scala 348:39]
  wire  _T_879 = _T_872 & _T_875; // @[GraphicEngineVGA.scala 350:59]
  wire  _T_880 = _T_879 & _T_878; // @[GraphicEngineVGA.scala 350:72]
  wire  _T_881 = _T_875 & _T_878; // @[GraphicEngineVGA.scala 350:97]
  wire [6:0] _T_892 = {{2'd0}, inSpriteX_6[4:0]}; // @[Mux.scala 80:57]
  wire [6:0] _T_904 = {{2'd0}, inSpriteY_6[4:0]}; // @[Mux.scala 80:57]
  wire [12:0] _T_907 = 7'h20 * _T_904; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_68021 = {{6'd0}, _T_892}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_909 = _GEN_68021 + _T_907; // @[GraphicEngineVGA.scala 367:46]
  wire [11:0] _T_912 = $signed(_T_232) - 11'sh0; // @[GraphicEngineVGA.scala 301:73]
  wire [11:0] _T_922 = $signed(_T_242) - 11'sh0; // @[GraphicEngineVGA.scala 302:73]
  wire [10:0] inSpriteY_7 = _T_922[10:0]; // @[GraphicEngineVGA.scala 263:23 GraphicEngineVGA.scala 322:18]
  wire  _T_963 = $signed(_T_912) >= 12'sh0; // @[GraphicEngineVGA.scala 343:27]
  wire  _T_971 = $signed(_T_912) < 12'sh20; // @[GraphicEngineVGA.scala 347:52]
  wire  _T_972 = _T_963 & _T_971; // @[GraphicEngineVGA.scala 347:39]
  wire  _T_973 = $signed(inSpriteY_7) >= 11'sh0; // @[GraphicEngineVGA.scala 348:31]
  wire  _T_974 = $signed(inSpriteY_7) < 11'sh20; // @[GraphicEngineVGA.scala 348:52]
  wire  _T_975 = _T_973 & _T_974; // @[GraphicEngineVGA.scala 348:39]
  wire [6:0] _T_989 = {{2'd0}, _T_912[4:0]}; // @[Mux.scala 80:57]
  wire [6:0] _T_1001 = {{2'd0}, inSpriteY_7[4:0]}; // @[Mux.scala 80:57]
  wire [12:0] _T_1004 = 7'h20 * _T_1001; // @[GraphicEngineVGA.scala 367:58]
  wire [12:0] _GEN_68026 = {{6'd0}, _T_989}; // @[GraphicEngineVGA.scala 367:46]
  wire [12:0] _T_1006 = _GEN_68026 + _T_1004; // @[GraphicEngineVGA.scala 367:46]
  reg [5:0] _T_1784; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1786_0; // @[GameUtilities.scala 21:24]
  reg  _T_1786_1; // @[GameUtilities.scala 21:24]
  reg  _T_1789; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1790 = ~_T_1789; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1793; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1795_0; // @[GameUtilities.scala 21:24]
  reg  _T_1795_1; // @[GameUtilities.scala 21:24]
  reg  _T_1798; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1799 = ~_T_1798; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1802; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1804_0; // @[GameUtilities.scala 21:24]
  reg  _T_1804_1; // @[GameUtilities.scala 21:24]
  reg  _T_1807; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1808 = ~_T_1807; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1811; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1813_0; // @[GameUtilities.scala 21:24]
  reg  _T_1813_1; // @[GameUtilities.scala 21:24]
  reg  _T_1816; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1817 = ~_T_1816; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1820; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1822_0; // @[GameUtilities.scala 21:24]
  reg  _T_1822_1; // @[GameUtilities.scala 21:24]
  reg  _T_1825; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1826 = ~_T_1825; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1829; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1831_0; // @[GameUtilities.scala 21:24]
  reg  _T_1831_1; // @[GameUtilities.scala 21:24]
  reg  _T_1834; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1835 = ~_T_1834; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1838; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1840_0; // @[GameUtilities.scala 21:24]
  reg  _T_1840_1; // @[GameUtilities.scala 21:24]
  reg  _T_1843; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1844 = ~_T_1843; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1847; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1848_0; // @[GameUtilities.scala 21:24]
  reg  _T_1848_1; // @[GameUtilities.scala 21:24]
  reg  _T_1849_0; // @[GameUtilities.scala 21:24]
  reg  _T_1849_1; // @[GameUtilities.scala 21:24]
  wire  _T_1850 = _T_1848_0 & _T_1849_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1852; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1853 = ~_T_1852; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1856; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1857_0; // @[GameUtilities.scala 21:24]
  reg  _T_1857_1; // @[GameUtilities.scala 21:24]
  reg  _T_1858_0; // @[GameUtilities.scala 21:24]
  reg  _T_1858_1; // @[GameUtilities.scala 21:24]
  wire  _T_1859 = _T_1857_0 & _T_1858_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1861; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1862 = ~_T_1861; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1865; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1866_0; // @[GameUtilities.scala 21:24]
  reg  _T_1866_1; // @[GameUtilities.scala 21:24]
  reg  _T_1867_0; // @[GameUtilities.scala 21:24]
  reg  _T_1867_1; // @[GameUtilities.scala 21:24]
  wire  _T_1868 = _T_1866_0 & _T_1867_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1870; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1871 = ~_T_1870; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1874; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1875_0; // @[GameUtilities.scala 21:24]
  reg  _T_1875_1; // @[GameUtilities.scala 21:24]
  reg  _T_1876_0; // @[GameUtilities.scala 21:24]
  reg  _T_1876_1; // @[GameUtilities.scala 21:24]
  wire  _T_1877 = _T_1875_0 & _T_1876_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1879; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1880 = ~_T_1879; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1883; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1884_0; // @[GameUtilities.scala 21:24]
  reg  _T_1884_1; // @[GameUtilities.scala 21:24]
  reg  _T_1885_0; // @[GameUtilities.scala 21:24]
  reg  _T_1885_1; // @[GameUtilities.scala 21:24]
  wire  _T_1886 = _T_1884_0 & _T_1885_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1888; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1889 = ~_T_1888; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1892; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1893_0; // @[GameUtilities.scala 21:24]
  reg  _T_1893_1; // @[GameUtilities.scala 21:24]
  reg  _T_1894_0; // @[GameUtilities.scala 21:24]
  reg  _T_1894_1; // @[GameUtilities.scala 21:24]
  wire  _T_1895 = _T_1893_0 & _T_1894_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1897; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1898 = ~_T_1897; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1901; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1902_0; // @[GameUtilities.scala 21:24]
  reg  _T_1902_1; // @[GameUtilities.scala 21:24]
  reg  _T_1903_0; // @[GameUtilities.scala 21:24]
  reg  _T_1903_1; // @[GameUtilities.scala 21:24]
  wire  _T_1904 = _T_1902_0 & _T_1903_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1906; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1907 = ~_T_1906; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1910; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1911_0; // @[GameUtilities.scala 21:24]
  reg  _T_1911_1; // @[GameUtilities.scala 21:24]
  reg  _T_1912_0; // @[GameUtilities.scala 21:24]
  reg  _T_1912_1; // @[GameUtilities.scala 21:24]
  wire  _T_1913 = _T_1911_0 & _T_1912_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1915; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1916 = ~_T_1915; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] _T_1919; // @[GraphicEngineVGA.scala 374:60]
  reg  _T_1920_0; // @[GameUtilities.scala 21:24]
  reg  _T_1920_1; // @[GameUtilities.scala 21:24]
  reg  _T_1921_0; // @[GameUtilities.scala 21:24]
  reg  _T_1921_1; // @[GameUtilities.scala 21:24]
  wire  _T_1922 = _T_1920_0 & _T_1921_0; // @[GraphicEngineVGA.scala 375:91]
  reg  _T_1924; // @[GraphicEngineVGA.scala 375:132]
  wire  _T_1925 = ~_T_1924; // @[GraphicEngineVGA.scala 375:123]
  reg [5:0] pixelColorSprite; // @[GraphicEngineVGA.scala 377:33]
  reg  pixelColorSpriteValid; // @[GraphicEngineVGA.scala 378:38]
  wire [5:0] pixelColorInDisplay = pixelColorSpriteValid ? pixelColorSprite : pixelColorBack; // @[GraphicEngineVGA.scala 382:32]
  reg  _T_1927_0; // @[GameUtilities.scala 21:24]
  reg  _T_1927_1; // @[GameUtilities.scala 21:24]
  reg  _T_1927_2; // @[GameUtilities.scala 21:24]
  wire [5:0] pixelColourVGA = _T_1927_0 ? pixelColorInDisplay : 6'h0; // @[GraphicEngineVGA.scala 383:27]
  reg [3:0] _T_1934; // @[GraphicEngineVGA.scala 387:23]
  reg [3:0] _T_1935; // @[GraphicEngineVGA.scala 388:25]
  reg [3:0] _T_1936; // @[GraphicEngineVGA.scala 389:24]
  Memory backTileMemories_0 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_0_clock),
    .io_address(backTileMemories_0_io_address),
    .io_dataRead(backTileMemories_0_io_dataRead)
  );
  Memory_1 backTileMemories_1 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_1_clock),
    .io_address(backTileMemories_1_io_address),
    .io_dataRead(backTileMemories_1_io_dataRead)
  );
  Memory_2 backTileMemories_2 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_2_clock),
    .io_address(backTileMemories_2_io_address),
    .io_dataRead(backTileMemories_2_io_dataRead)
  );
  Memory_3 backTileMemories_3 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_3_clock),
    .io_address(backTileMemories_3_io_address),
    .io_dataRead(backTileMemories_3_io_dataRead)
  );
  Memory_4 backTileMemories_4 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_4_clock),
    .io_address(backTileMemories_4_io_address),
    .io_dataRead(backTileMemories_4_io_dataRead)
  );
  Memory_5 backTileMemories_5 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_5_clock),
    .io_address(backTileMemories_5_io_address),
    .io_dataRead(backTileMemories_5_io_dataRead)
  );
  Memory_6 backTileMemories_6 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_6_clock),
    .io_address(backTileMemories_6_io_address),
    .io_dataRead(backTileMemories_6_io_dataRead)
  );
  Memory_7 backTileMemories_7 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_7_clock),
    .io_address(backTileMemories_7_io_address),
    .io_dataRead(backTileMemories_7_io_dataRead)
  );
  Memory_8 backTileMemories_8 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_8_clock),
    .io_address(backTileMemories_8_io_address),
    .io_dataRead(backTileMemories_8_io_dataRead)
  );
  Memory_9 backTileMemories_9 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_9_clock),
    .io_address(backTileMemories_9_io_address),
    .io_dataRead(backTileMemories_9_io_dataRead)
  );
  Memory_10 backTileMemories_10 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_10_clock),
    .io_address(backTileMemories_10_io_address),
    .io_dataRead(backTileMemories_10_io_dataRead)
  );
  Memory_11 backTileMemories_11 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_11_clock),
    .io_address(backTileMemories_11_io_address),
    .io_dataRead(backTileMemories_11_io_dataRead)
  );
  Memory_12 backTileMemories_12 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_12_clock),
    .io_address(backTileMemories_12_io_address),
    .io_dataRead(backTileMemories_12_io_dataRead)
  );
  Memory_13 backTileMemories_13 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_13_clock),
    .io_address(backTileMemories_13_io_address),
    .io_dataRead(backTileMemories_13_io_dataRead)
  );
  Memory_14 backTileMemories_14 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_14_clock),
    .io_address(backTileMemories_14_io_address),
    .io_dataRead(backTileMemories_14_io_dataRead)
  );
  Memory_15 backTileMemories_15 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_15_clock),
    .io_address(backTileMemories_15_io_address),
    .io_dataRead(backTileMemories_15_io_dataRead)
  );
  Memory_16 backTileMemories_16 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_16_clock),
    .io_address(backTileMemories_16_io_address),
    .io_dataRead(backTileMemories_16_io_dataRead)
  );
  Memory_17 backTileMemories_17 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_17_clock),
    .io_address(backTileMemories_17_io_address),
    .io_dataRead(backTileMemories_17_io_dataRead)
  );
  Memory_18 backTileMemories_18 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_18_clock),
    .io_address(backTileMemories_18_io_address),
    .io_dataRead(backTileMemories_18_io_dataRead)
  );
  Memory_19 backTileMemories_19 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_19_clock),
    .io_address(backTileMemories_19_io_address),
    .io_dataRead(backTileMemories_19_io_dataRead)
  );
  Memory_20 backTileMemories_20 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_20_clock),
    .io_address(backTileMemories_20_io_address),
    .io_dataRead(backTileMemories_20_io_dataRead)
  );
  Memory_21 backTileMemories_21 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_21_clock),
    .io_address(backTileMemories_21_io_address),
    .io_dataRead(backTileMemories_21_io_dataRead)
  );
  Memory_22 backTileMemories_22 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_22_clock),
    .io_address(backTileMemories_22_io_address),
    .io_dataRead(backTileMemories_22_io_dataRead)
  );
  Memory_23 backTileMemories_23 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_23_clock),
    .io_address(backTileMemories_23_io_address),
    .io_dataRead(backTileMemories_23_io_dataRead)
  );
  Memory_24 backTileMemories_24 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_24_clock),
    .io_address(backTileMemories_24_io_address),
    .io_dataRead(backTileMemories_24_io_dataRead)
  );
  Memory_25 backTileMemories_25 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_25_clock),
    .io_address(backTileMemories_25_io_address),
    .io_dataRead(backTileMemories_25_io_dataRead)
  );
  Memory_26 backTileMemories_26 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_26_clock),
    .io_address(backTileMemories_26_io_address),
    .io_dataRead(backTileMemories_26_io_dataRead)
  );
  Memory_27 backTileMemories_27 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_27_clock),
    .io_address(backTileMemories_27_io_address),
    .io_dataRead(backTileMemories_27_io_dataRead)
  );
  Memory_28 backTileMemories_28 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_28_clock),
    .io_address(backTileMemories_28_io_address),
    .io_dataRead(backTileMemories_28_io_dataRead)
  );
  Memory_29 backTileMemories_29 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_29_clock),
    .io_address(backTileMemories_29_io_address),
    .io_dataRead(backTileMemories_29_io_dataRead)
  );
  Memory_30 backTileMemories_30 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_30_clock),
    .io_address(backTileMemories_30_io_address),
    .io_dataRead(backTileMemories_30_io_dataRead)
  );
  Memory_31 backTileMemories_31 ( // @[GraphicEngineVGA.scala 165:32]
    .clock(backTileMemories_31_clock),
    .io_address(backTileMemories_31_io_address),
    .io_dataRead(backTileMemories_31_io_dataRead)
  );
  Memory_32 backBufferMemory ( // @[GraphicEngineVGA.scala 182:32]
    .clock(backBufferMemory_clock),
    .io_address(backBufferMemory_io_address),
    .io_dataRead(backBufferMemory_io_dataRead),
    .io_writeEnable(backBufferMemory_io_writeEnable),
    .io_dataWrite(backBufferMemory_io_dataWrite)
  );
  Memory_32 backBufferShadowMemory ( // @[GraphicEngineVGA.scala 183:38]
    .clock(backBufferShadowMemory_clock),
    .io_address(backBufferShadowMemory_io_address),
    .io_dataRead(backBufferShadowMemory_io_dataRead),
    .io_writeEnable(backBufferShadowMemory_io_writeEnable),
    .io_dataWrite(backBufferShadowMemory_io_dataWrite)
  );
  Memory_34 backBufferRestoreMemory ( // @[GraphicEngineVGA.scala 184:39]
    .clock(backBufferRestoreMemory_clock),
    .io_address(backBufferRestoreMemory_io_address),
    .io_dataRead(backBufferRestoreMemory_io_dataRead)
  );
  Memory_35 spriteMemories_0 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_0_clock),
    .io_address(spriteMemories_0_io_address),
    .io_dataRead(spriteMemories_0_io_dataRead)
  );
  Memory_36 spriteMemories_1 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_1_clock),
    .io_address(spriteMemories_1_io_address),
    .io_dataRead(spriteMemories_1_io_dataRead)
  );
  Memory_37 spriteMemories_2 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_2_clock),
    .io_address(spriteMemories_2_io_address),
    .io_dataRead(spriteMemories_2_io_dataRead)
  );
  Memory_38 spriteMemories_3 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_3_clock),
    .io_address(spriteMemories_3_io_address),
    .io_dataRead(spriteMemories_3_io_dataRead)
  );
  Memory_39 spriteMemories_4 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_4_clock),
    .io_address(spriteMemories_4_io_address),
    .io_dataRead(spriteMemories_4_io_dataRead)
  );
  Memory_40 spriteMemories_5 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_5_clock),
    .io_address(spriteMemories_5_io_address),
    .io_dataRead(spriteMemories_5_io_dataRead)
  );
  Memory_41 spriteMemories_6 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_6_clock),
    .io_address(spriteMemories_6_io_address),
    .io_dataRead(spriteMemories_6_io_dataRead)
  );
  Memory_42 spriteMemories_7 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_7_clock),
    .io_address(spriteMemories_7_io_address),
    .io_dataRead(spriteMemories_7_io_dataRead)
  );
  Memory_43 spriteMemories_8 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_8_clock),
    .io_address(spriteMemories_8_io_address),
    .io_dataRead(spriteMemories_8_io_dataRead)
  );
  Memory_44 spriteMemories_9 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_9_clock),
    .io_address(spriteMemories_9_io_address),
    .io_dataRead(spriteMemories_9_io_dataRead)
  );
  Memory_45 spriteMemories_10 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_10_clock),
    .io_address(spriteMemories_10_io_address),
    .io_dataRead(spriteMemories_10_io_dataRead)
  );
  Memory_46 spriteMemories_11 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_11_clock),
    .io_address(spriteMemories_11_io_address),
    .io_dataRead(spriteMemories_11_io_dataRead)
  );
  Memory_47 spriteMemories_12 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_12_clock),
    .io_address(spriteMemories_12_io_address),
    .io_dataRead(spriteMemories_12_io_dataRead)
  );
  Memory_48 spriteMemories_13 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_13_clock),
    .io_address(spriteMemories_13_io_address),
    .io_dataRead(spriteMemories_13_io_dataRead)
  );
  Memory_49 spriteMemories_14 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_14_clock),
    .io_address(spriteMemories_14_io_address),
    .io_dataRead(spriteMemories_14_io_dataRead)
  );
  Memory_50 spriteMemories_15 ( // @[GraphicEngineVGA.scala 254:30]
    .clock(spriteMemories_15_clock),
    .io_address(spriteMemories_15_io_address),
    .io_dataRead(spriteMemories_15_io_dataRead)
  );
  MultiHotPriortyReductionTree multiHotPriortyReductionTree ( // @[GraphicEngineVGA.scala 372:44]
    .io_dataInput_0(multiHotPriortyReductionTree_io_dataInput_0),
    .io_dataInput_1(multiHotPriortyReductionTree_io_dataInput_1),
    .io_dataInput_2(multiHotPriortyReductionTree_io_dataInput_2),
    .io_dataInput_3(multiHotPriortyReductionTree_io_dataInput_3),
    .io_dataInput_4(multiHotPriortyReductionTree_io_dataInput_4),
    .io_dataInput_5(multiHotPriortyReductionTree_io_dataInput_5),
    .io_dataInput_6(multiHotPriortyReductionTree_io_dataInput_6),
    .io_dataInput_7(multiHotPriortyReductionTree_io_dataInput_7),
    .io_dataInput_8(multiHotPriortyReductionTree_io_dataInput_8),
    .io_dataInput_9(multiHotPriortyReductionTree_io_dataInput_9),
    .io_dataInput_10(multiHotPriortyReductionTree_io_dataInput_10),
    .io_dataInput_11(multiHotPriortyReductionTree_io_dataInput_11),
    .io_dataInput_12(multiHotPriortyReductionTree_io_dataInput_12),
    .io_dataInput_13(multiHotPriortyReductionTree_io_dataInput_13),
    .io_dataInput_14(multiHotPriortyReductionTree_io_dataInput_14),
    .io_dataInput_15(multiHotPriortyReductionTree_io_dataInput_15),
    .io_selectInput_0(multiHotPriortyReductionTree_io_selectInput_0),
    .io_selectInput_1(multiHotPriortyReductionTree_io_selectInput_1),
    .io_selectInput_2(multiHotPriortyReductionTree_io_selectInput_2),
    .io_selectInput_3(multiHotPriortyReductionTree_io_selectInput_3),
    .io_selectInput_4(multiHotPriortyReductionTree_io_selectInput_4),
    .io_selectInput_5(multiHotPriortyReductionTree_io_selectInput_5),
    .io_selectInput_6(multiHotPriortyReductionTree_io_selectInput_6),
    .io_selectInput_7(multiHotPriortyReductionTree_io_selectInput_7),
    .io_selectInput_8(multiHotPriortyReductionTree_io_selectInput_8),
    .io_selectInput_9(multiHotPriortyReductionTree_io_selectInput_9),
    .io_selectInput_10(multiHotPriortyReductionTree_io_selectInput_10),
    .io_selectInput_11(multiHotPriortyReductionTree_io_selectInput_11),
    .io_selectInput_12(multiHotPriortyReductionTree_io_selectInput_12),
    .io_selectInput_13(multiHotPriortyReductionTree_io_selectInput_13),
    .io_selectInput_14(multiHotPriortyReductionTree_io_selectInput_14),
    .io_selectInput_15(multiHotPriortyReductionTree_io_selectInput_15),
    .io_dataOutput(multiHotPriortyReductionTree_io_dataOutput),
    .io_selectOutput(multiHotPriortyReductionTree_io_selectOutput)
  );
  assign io_newFrame = run & _GEN_8; // @[GraphicEngineVGA.scala 73:15 GraphicEngineVGA.scala 83:23]
  assign io_missingFrameError = missingFrameErrorReg; // @[GraphicEngineVGA.scala 135:24]
  assign io_vgaRed = _T_1934; // @[GraphicEngineVGA.scala 387:13]
  assign io_vgaBlue = _T_1936; // @[GraphicEngineVGA.scala 389:14]
  assign io_vgaGreen = _T_1935; // @[GraphicEngineVGA.scala 388:15]
  assign io_Hsync = _T_14_0; // @[GraphicEngineVGA.scala 97:12]
  assign io_Vsync = _T_16_0; // @[GraphicEngineVGA.scala 98:12]
  assign backTileMemories_0_clock = clock;
  assign backTileMemories_0_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_1_clock = clock;
  assign backTileMemories_1_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_2_clock = clock;
  assign backTileMemories_2_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_3_clock = clock;
  assign backTileMemories_3_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_4_clock = clock;
  assign backTileMemories_4_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_5_clock = clock;
  assign backTileMemories_5_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_6_clock = clock;
  assign backTileMemories_6_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_7_clock = clock;
  assign backTileMemories_7_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_8_clock = clock;
  assign backTileMemories_8_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_9_clock = clock;
  assign backTileMemories_9_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_10_clock = clock;
  assign backTileMemories_10_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_11_clock = clock;
  assign backTileMemories_11_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_12_clock = clock;
  assign backTileMemories_12_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_13_clock = clock;
  assign backTileMemories_13_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_14_clock = clock;
  assign backTileMemories_14_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_15_clock = clock;
  assign backTileMemories_15_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_16_clock = clock;
  assign backTileMemories_16_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_17_clock = clock;
  assign backTileMemories_17_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_18_clock = clock;
  assign backTileMemories_18_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_19_clock = clock;
  assign backTileMemories_19_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_20_clock = clock;
  assign backTileMemories_20_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_21_clock = clock;
  assign backTileMemories_21_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_22_clock = clock;
  assign backTileMemories_22_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_23_clock = clock;
  assign backTileMemories_23_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_24_clock = clock;
  assign backTileMemories_24_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_25_clock = clock;
  assign backTileMemories_25_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_26_clock = clock;
  assign backTileMemories_26_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_27_clock = clock;
  assign backTileMemories_27_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_28_clock = clock;
  assign backTileMemories_28_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_29_clock = clock;
  assign backTileMemories_29_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_30_clock = clock;
  assign backTileMemories_30_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backTileMemories_31_clock = clock;
  assign backTileMemories_31_io_address = _T_41[9:0]; // @[GraphicEngineVGA.scala 176:36]
  assign backBufferMemory_clock = clock;
  assign backBufferMemory_io_address = _T_223[10:0]; // @[GraphicEngineVGA.scala 230:31]
  assign backBufferMemory_io_writeEnable = copyEnabledReg; // @[GraphicEngineVGA.scala 232:35]
  assign backBufferMemory_io_dataWrite = backBufferShadowMemory_io_dataRead; // @[GraphicEngineVGA.scala 233:33]
  assign backBufferShadowMemory_clock = clock;
  assign backBufferShadowMemory_io_address = restoreEnabled ? _T_206 : _T_209; // @[GraphicEngineVGA.scala 225:37]
  assign backBufferShadowMemory_io_writeEnable = restoreEnabled & _T_211; // @[GraphicEngineVGA.scala 227:41]
  assign backBufferShadowMemory_io_dataWrite = restoreEnabled ? backBufferRestoreMemory_io_dataRead : 5'h0; // @[GraphicEngineVGA.scala 228:39]
  assign backBufferRestoreMemory_clock = clock;
  assign backBufferRestoreMemory_io_address = backMemoryRestoreCounter[10:0]; // @[GraphicEngineVGA.scala 220:38]
  assign spriteMemories_0_clock = clock;
  assign spriteMemories_0_io_address = _T_327[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_1_clock = clock;
  assign spriteMemories_1_io_address = _T_424[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_2_clock = clock;
  assign spriteMemories_2_io_address = _T_521[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_3_clock = clock;
  assign spriteMemories_3_io_address = _T_618[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_4_clock = clock;
  assign spriteMemories_4_io_address = _T_715[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_5_clock = clock;
  assign spriteMemories_5_io_address = _T_812[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_6_clock = clock;
  assign spriteMemories_6_io_address = _T_909[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_7_clock = clock;
  assign spriteMemories_7_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_8_clock = clock;
  assign spriteMemories_8_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_9_clock = clock;
  assign spriteMemories_9_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_10_clock = clock;
  assign spriteMemories_10_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_11_clock = clock;
  assign spriteMemories_11_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_12_clock = clock;
  assign spriteMemories_12_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_13_clock = clock;
  assign spriteMemories_13_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_14_clock = clock;
  assign spriteMemories_14_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign spriteMemories_15_clock = clock;
  assign spriteMemories_15_io_address = _T_1006[9:0]; // @[GraphicEngineVGA.scala 367:38]
  assign multiHotPriortyReductionTree_io_dataInput_0 = _T_1784; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_1 = _T_1793; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_2 = _T_1802; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_3 = _T_1811; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_4 = _T_1820; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_5 = _T_1829; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_6 = _T_1838; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_7 = _T_1847; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_8 = _T_1856; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_9 = _T_1865; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_10 = _T_1874; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_11 = _T_1883; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_12 = _T_1892; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_13 = _T_1901; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_14 = _T_1910; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_dataInput_15 = _T_1919; // @[GraphicEngineVGA.scala 374:50]
  assign multiHotPriortyReductionTree_io_selectInput_0 = _T_1786_0 & _T_1790; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_1 = _T_1795_0 & _T_1799; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_2 = _T_1804_0 & _T_1808; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_3 = _T_1813_0 & _T_1817; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_4 = _T_1822_0 & _T_1826; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_5 = _T_1831_0 & _T_1835; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_6 = _T_1840_0 & _T_1844; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_7 = _T_1850 & _T_1853; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_8 = _T_1859 & _T_1862; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_9 = _T_1868 & _T_1871; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_10 = _T_1877 & _T_1880; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_11 = _T_1886 & _T_1889; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_12 = _T_1895 & _T_1898; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_13 = _T_1904 & _T_1907; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_14 = _T_1913 & _T_1916; // @[GraphicEngineVGA.scala 375:52]
  assign multiHotPriortyReductionTree_io_selectInput_15 = _T_1922 & _T_1925; // @[GraphicEngineVGA.scala 375:52]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ScaleCounterReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  CounterXReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  CounterYReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  backMemoryRestoreCounter = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  _T_14_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_14_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_14_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_14_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_16_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_16_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_16_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_16_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  frameClockCount = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXPositionReg_0 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXPositionReg_1 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXPositionReg_2 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXPositionReg_3 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXPositionReg_4 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXPositionReg_5 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXPositionReg_6 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteYPositionReg_0 = _RAND_20[9:0];
  _RAND_21 = {1{`RANDOM}};
  spriteYPositionReg_1 = _RAND_21[9:0];
  _RAND_22 = {1{`RANDOM}};
  spriteYPositionReg_2 = _RAND_22[9:0];
  _RAND_23 = {1{`RANDOM}};
  spriteYPositionReg_3 = _RAND_23[9:0];
  _RAND_24 = {1{`RANDOM}};
  spriteYPositionReg_4 = _RAND_24[9:0];
  _RAND_25 = {1{`RANDOM}};
  spriteYPositionReg_5 = _RAND_25[9:0];
  _RAND_26 = {1{`RANDOM}};
  spriteYPositionReg_6 = _RAND_26[9:0];
  _RAND_27 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  spriteFlipHorizontalReg_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  spriteFlipHorizontalReg_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  spriteFlipHorizontalReg_4 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  spriteFlipVerticalReg_2 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  spriteFlipVerticalReg_5 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  spriteScaleHorizontalReg_0 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  spriteScaleHorizontalReg_1 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  spriteScaleHorizontalReg_2 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  spriteScaleHorizontalReg_4 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  spriteScaleVerticalReg_0 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  spriteScaleVerticalReg_1 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  spriteScaleVerticalReg_2 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  spriteScaleVerticalReg_4 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  spriteRotationReg_4 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  spriteRotationReg_6 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  missingFrameErrorReg = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  newFrameStikyReg = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_36 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  backTileMemoryDataRead_0 = _RAND_54[6:0];
  _RAND_55 = {1{`RANDOM}};
  backTileMemoryDataRead_1 = _RAND_55[6:0];
  _RAND_56 = {1{`RANDOM}};
  backTileMemoryDataRead_2 = _RAND_56[6:0];
  _RAND_57 = {1{`RANDOM}};
  backTileMemoryDataRead_3 = _RAND_57[6:0];
  _RAND_58 = {1{`RANDOM}};
  backTileMemoryDataRead_4 = _RAND_58[6:0];
  _RAND_59 = {1{`RANDOM}};
  backTileMemoryDataRead_5 = _RAND_59[6:0];
  _RAND_60 = {1{`RANDOM}};
  backTileMemoryDataRead_6 = _RAND_60[6:0];
  _RAND_61 = {1{`RANDOM}};
  backTileMemoryDataRead_7 = _RAND_61[6:0];
  _RAND_62 = {1{`RANDOM}};
  backTileMemoryDataRead_8 = _RAND_62[6:0];
  _RAND_63 = {1{`RANDOM}};
  backTileMemoryDataRead_9 = _RAND_63[6:0];
  _RAND_64 = {1{`RANDOM}};
  backTileMemoryDataRead_10 = _RAND_64[6:0];
  _RAND_65 = {1{`RANDOM}};
  backTileMemoryDataRead_11 = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  backTileMemoryDataRead_12 = _RAND_66[6:0];
  _RAND_67 = {1{`RANDOM}};
  backTileMemoryDataRead_13 = _RAND_67[6:0];
  _RAND_68 = {1{`RANDOM}};
  backTileMemoryDataRead_14 = _RAND_68[6:0];
  _RAND_69 = {1{`RANDOM}};
  backTileMemoryDataRead_15 = _RAND_69[6:0];
  _RAND_70 = {1{`RANDOM}};
  backTileMemoryDataRead_16 = _RAND_70[6:0];
  _RAND_71 = {1{`RANDOM}};
  backTileMemoryDataRead_17 = _RAND_71[6:0];
  _RAND_72 = {1{`RANDOM}};
  backTileMemoryDataRead_18 = _RAND_72[6:0];
  _RAND_73 = {1{`RANDOM}};
  backTileMemoryDataRead_19 = _RAND_73[6:0];
  _RAND_74 = {1{`RANDOM}};
  backTileMemoryDataRead_20 = _RAND_74[6:0];
  _RAND_75 = {1{`RANDOM}};
  backTileMemoryDataRead_21 = _RAND_75[6:0];
  _RAND_76 = {1{`RANDOM}};
  backTileMemoryDataRead_22 = _RAND_76[6:0];
  _RAND_77 = {1{`RANDOM}};
  backTileMemoryDataRead_23 = _RAND_77[6:0];
  _RAND_78 = {1{`RANDOM}};
  backTileMemoryDataRead_24 = _RAND_78[6:0];
  _RAND_79 = {1{`RANDOM}};
  backTileMemoryDataRead_25 = _RAND_79[6:0];
  _RAND_80 = {1{`RANDOM}};
  backTileMemoryDataRead_26 = _RAND_80[6:0];
  _RAND_81 = {1{`RANDOM}};
  backTileMemoryDataRead_27 = _RAND_81[6:0];
  _RAND_82 = {1{`RANDOM}};
  backTileMemoryDataRead_28 = _RAND_82[6:0];
  _RAND_83 = {1{`RANDOM}};
  backTileMemoryDataRead_29 = _RAND_83[6:0];
  _RAND_84 = {1{`RANDOM}};
  backTileMemoryDataRead_30 = _RAND_84[6:0];
  _RAND_85 = {1{`RANDOM}};
  backTileMemoryDataRead_31 = _RAND_85[6:0];
  _RAND_86 = {1{`RANDOM}};
  backMemoryCopyCounter = _RAND_86[11:0];
  _RAND_87 = {1{`RANDOM}};
  copyEnabledReg = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _T_206 = _RAND_88[10:0];
  _RAND_89 = {1{`RANDOM}};
  _T_211 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _T_218 = _RAND_90[10:0];
  _RAND_91 = {1{`RANDOM}};
  _T_225 = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  pixelColorBack = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  _T_1784 = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  _T_1786_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _T_1786_1 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _T_1789 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _T_1793 = _RAND_97[5:0];
  _RAND_98 = {1{`RANDOM}};
  _T_1795_0 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _T_1795_1 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _T_1798 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  _T_1802 = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  _T_1804_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  _T_1804_1 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  _T_1807 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _T_1811 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  _T_1813_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  _T_1813_1 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _T_1816 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  _T_1820 = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  _T_1822_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  _T_1822_1 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  _T_1825 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  _T_1829 = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  _T_1831_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  _T_1831_1 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  _T_1834 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  _T_1838 = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  _T_1840_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  _T_1840_1 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  _T_1843 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  _T_1847 = _RAND_121[5:0];
  _RAND_122 = {1{`RANDOM}};
  _T_1848_0 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  _T_1848_1 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  _T_1849_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  _T_1849_1 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  _T_1852 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  _T_1856 = _RAND_127[5:0];
  _RAND_128 = {1{`RANDOM}};
  _T_1857_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  _T_1857_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  _T_1858_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  _T_1858_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  _T_1861 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _T_1865 = _RAND_133[5:0];
  _RAND_134 = {1{`RANDOM}};
  _T_1866_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  _T_1866_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _T_1867_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  _T_1867_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _T_1870 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  _T_1874 = _RAND_139[5:0];
  _RAND_140 = {1{`RANDOM}};
  _T_1875_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  _T_1875_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _T_1876_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  _T_1876_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _T_1879 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  _T_1883 = _RAND_145[5:0];
  _RAND_146 = {1{`RANDOM}};
  _T_1884_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _T_1884_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _T_1885_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  _T_1885_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _T_1888 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  _T_1892 = _RAND_151[5:0];
  _RAND_152 = {1{`RANDOM}};
  _T_1893_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  _T_1893_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _T_1894_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  _T_1894_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _T_1897 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _T_1901 = _RAND_157[5:0];
  _RAND_158 = {1{`RANDOM}};
  _T_1902_0 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  _T_1902_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _T_1903_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  _T_1903_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _T_1906 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  _T_1910 = _RAND_163[5:0];
  _RAND_164 = {1{`RANDOM}};
  _T_1911_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _T_1911_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _T_1912_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_1912_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  _T_1915 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  _T_1919 = _RAND_169[5:0];
  _RAND_170 = {1{`RANDOM}};
  _T_1920_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  _T_1920_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _T_1921_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  _T_1921_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_1924 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  pixelColorSprite = _RAND_175[5:0];
  _RAND_176 = {1{`RANDOM}};
  pixelColorSpriteValid = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_1927_0 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _T_1927_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _T_1927_2 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _T_1934 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  _T_1935 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  _T_1936 = _RAND_182[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ScaleCounterReg <= 2'h0;
    end else if (run) begin
      if (_T) begin
        ScaleCounterReg <= 2'h0;
      end else begin
        ScaleCounterReg <= _T_8;
      end
    end
    if (reset) begin
      CounterXReg <= 10'h0;
    end else if (run) begin
      if (_T) begin
        if (_T_1) begin
          CounterXReg <= 10'h0;
        end else begin
          CounterXReg <= _T_6;
        end
      end
    end
    if (reset) begin
      CounterYReg <= 10'h0;
    end else if (run) begin
      if (_T) begin
        if (_T_1) begin
          if (_T_2) begin
            CounterYReg <= 10'h0;
          end else begin
            CounterYReg <= _T_4;
          end
        end
      end
    end
    if (reset) begin
      backMemoryRestoreCounter <= 12'h0;
    end else if (restoreEnabled) begin
      backMemoryRestoreCounter <= _T_203;
    end
    _T_14_0 <= _T_14_1;
    _T_14_1 <= _T_14_2;
    _T_14_2 <= _T_14_3;
    _T_14_3 <= ~Hsync;
    _T_16_0 <= _T_16_1;
    _T_16_1 <= _T_16_2;
    _T_16_2 <= _T_16_3;
    _T_16_3 <= ~Vsync;
    if (reset) begin
      frameClockCount <= 21'h0;
    end else if (_T_19) begin
      frameClockCount <= 21'h0;
    end else begin
      frameClockCount <= _T_21;
    end
    if (reset) begin
      spriteXPositionReg_0 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_0 <= io_spriteXPosition_0;
    end
    if (reset) begin
      spriteXPositionReg_1 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_1 <= 11'sh96;
    end
    if (reset) begin
      spriteXPositionReg_2 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_2 <= 11'sh96;
    end
    if (reset) begin
      spriteXPositionReg_3 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_3 <= 11'sh96;
    end
    if (reset) begin
      spriteXPositionReg_4 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_4 <= 11'sh12c;
    end
    if (reset) begin
      spriteXPositionReg_5 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_5 <= 11'sh12c;
    end
    if (reset) begin
      spriteXPositionReg_6 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_6 <= 11'sh12c;
    end
    if (reset) begin
      spriteYPositionReg_0 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_0 <= io_spriteYPosition_0;
    end
    if (reset) begin
      spriteYPositionReg_1 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_1 <= 10'sh148;
    end
    if (reset) begin
      spriteYPositionReg_2 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_2 <= 10'sh148;
    end
    if (reset) begin
      spriteYPositionReg_3 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_3 <= 10'sh148;
    end
    if (reset) begin
      spriteYPositionReg_4 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_4 <= 10'sh148;
    end
    if (reset) begin
      spriteYPositionReg_5 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_5 <= 10'sh148;
    end
    if (reset) begin
      spriteYPositionReg_6 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_6 <= 10'sh148;
    end
    spriteVisibleReg_7 <= reset | _GEN_52;
    spriteVisibleReg_8 <= reset | _GEN_53;
    spriteVisibleReg_9 <= reset | _GEN_54;
    spriteVisibleReg_10 <= reset | _GEN_55;
    spriteVisibleReg_11 <= reset | _GEN_56;
    spriteVisibleReg_12 <= reset | _GEN_57;
    spriteVisibleReg_13 <= reset | _GEN_58;
    spriteVisibleReg_14 <= reset | _GEN_59;
    spriteVisibleReg_15 <= reset | _GEN_60;
    if (reset) begin
      spriteFlipHorizontalReg_0 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipHorizontalReg_0 <= io_spriteFlipHorizontal_0;
    end
    if (reset) begin
      spriteFlipHorizontalReg_1 <= 1'h0;
    end else begin
      spriteFlipHorizontalReg_1 <= _GEN_62;
    end
    if (reset) begin
      spriteFlipHorizontalReg_4 <= 1'h0;
    end else begin
      spriteFlipHorizontalReg_4 <= _GEN_65;
    end
    if (reset) begin
      spriteFlipVerticalReg_2 <= 1'h0;
    end else begin
      spriteFlipVerticalReg_2 <= _GEN_79;
    end
    if (reset) begin
      spriteFlipVerticalReg_5 <= 1'h0;
    end else begin
      spriteFlipVerticalReg_5 <= _GEN_82;
    end
    if (reset) begin
      spriteScaleHorizontalReg_0 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleHorizontalReg_0 <= 2'h1;
    end
    if (reset) begin
      spriteScaleHorizontalReg_1 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleHorizontalReg_1 <= 2'h1;
    end
    if (reset) begin
      spriteScaleHorizontalReg_2 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleHorizontalReg_2 <= 2'h1;
    end
    if (reset) begin
      spriteScaleHorizontalReg_4 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleHorizontalReg_4 <= 2'h1;
    end
    if (reset) begin
      spriteScaleVerticalReg_0 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleVerticalReg_0 <= 2'h2;
    end
    if (reset) begin
      spriteScaleVerticalReg_1 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleVerticalReg_1 <= 2'h1;
    end
    if (reset) begin
      spriteScaleVerticalReg_2 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleVerticalReg_2 <= 2'h1;
    end
    if (reset) begin
      spriteScaleVerticalReg_4 <= 2'h0;
    end else if (io_newFrame) begin
      spriteScaleVerticalReg_4 <= 2'h1;
    end
    if (reset) begin
      spriteRotationReg_4 <= 1'h0;
    end else begin
      spriteRotationReg_4 <= _GEN_129;
    end
    if (reset) begin
      spriteRotationReg_6 <= 1'h0;
    end else begin
      spriteRotationReg_6 <= _GEN_131;
    end
    if (reset) begin
      missingFrameErrorReg <= 1'h0;
    end else begin
      missingFrameErrorReg <= _GEN_146;
    end
    if (reset) begin
      newFrameStikyReg <= 1'h0;
    end else if (_T_36) begin
      newFrameStikyReg <= 1'h0;
    end else begin
      newFrameStikyReg <= _GEN_144;
    end
    _T_36 <= io_frameUpdateDone;
    backTileMemoryDataRead_0 <= backTileMemories_0_io_dataRead;
    backTileMemoryDataRead_1 <= backTileMemories_1_io_dataRead;
    backTileMemoryDataRead_2 <= backTileMemories_2_io_dataRead;
    backTileMemoryDataRead_3 <= backTileMemories_3_io_dataRead;
    backTileMemoryDataRead_4 <= backTileMemories_4_io_dataRead;
    backTileMemoryDataRead_5 <= backTileMemories_5_io_dataRead;
    backTileMemoryDataRead_6 <= backTileMemories_6_io_dataRead;
    backTileMemoryDataRead_7 <= backTileMemories_7_io_dataRead;
    backTileMemoryDataRead_8 <= backTileMemories_8_io_dataRead;
    backTileMemoryDataRead_9 <= backTileMemories_9_io_dataRead;
    backTileMemoryDataRead_10 <= backTileMemories_10_io_dataRead;
    backTileMemoryDataRead_11 <= backTileMemories_11_io_dataRead;
    backTileMemoryDataRead_12 <= backTileMemories_12_io_dataRead;
    backTileMemoryDataRead_13 <= backTileMemories_13_io_dataRead;
    backTileMemoryDataRead_14 <= backTileMemories_14_io_dataRead;
    backTileMemoryDataRead_15 <= backTileMemories_15_io_dataRead;
    backTileMemoryDataRead_16 <= backTileMemories_16_io_dataRead;
    backTileMemoryDataRead_17 <= backTileMemories_17_io_dataRead;
    backTileMemoryDataRead_18 <= backTileMemories_18_io_dataRead;
    backTileMemoryDataRead_19 <= backTileMemories_19_io_dataRead;
    backTileMemoryDataRead_20 <= backTileMemories_20_io_dataRead;
    backTileMemoryDataRead_21 <= backTileMemories_21_io_dataRead;
    backTileMemoryDataRead_22 <= backTileMemories_22_io_dataRead;
    backTileMemoryDataRead_23 <= backTileMemories_23_io_dataRead;
    backTileMemoryDataRead_24 <= backTileMemories_24_io_dataRead;
    backTileMemoryDataRead_25 <= backTileMemories_25_io_dataRead;
    backTileMemoryDataRead_26 <= backTileMemories_26_io_dataRead;
    backTileMemoryDataRead_27 <= backTileMemories_27_io_dataRead;
    backTileMemoryDataRead_28 <= backTileMemories_28_io_dataRead;
    backTileMemoryDataRead_29 <= backTileMemories_29_io_dataRead;
    backTileMemoryDataRead_30 <= backTileMemories_30_io_dataRead;
    backTileMemoryDataRead_31 <= backTileMemories_31_io_dataRead;
    if (reset) begin
      backMemoryCopyCounter <= 12'h0;
    end else if (preDisplayArea) begin
      if (_T_198) begin
        backMemoryCopyCounter <= _T_200;
      end
    end else begin
      backMemoryCopyCounter <= 12'h0;
    end
    copyEnabledReg <= preDisplayArea & _T_198;
    _T_206 <= backMemoryRestoreCounter[10:0];
    _T_211 <= backMemoryRestoreCounter < 12'h800;
    _T_218 <= backMemoryCopyCounter[10:0];
    _T_225 <= backBufferMemory_io_dataRead;
    if (fullBackgroundColor[6]) begin
      pixelColorBack <= 6'h0;
    end else begin
      pixelColorBack <= fullBackgroundColor[5:0];
    end
    _T_1784 <= spriteMemories_0_io_dataRead[5:0];
    _T_1786_0 <= _T_1786_1;
    _T_1786_1 <= _T_293 & _T_296;
    _T_1789 <= spriteMemories_0_io_dataRead[6];
    _T_1793 <= spriteMemories_1_io_dataRead[5:0];
    _T_1795_0 <= _T_1795_1;
    _T_1795_1 <= _T_390 & _T_393;
    _T_1798 <= spriteMemories_1_io_dataRead[6];
    _T_1802 <= spriteMemories_2_io_dataRead[5:0];
    _T_1804_0 <= _T_1804_1;
    _T_1804_1 <= _T_487 & _T_490;
    _T_1807 <= spriteMemories_2_io_dataRead[6];
    _T_1811 <= spriteMemories_3_io_dataRead[5:0];
    _T_1813_0 <= _T_1813_1;
    _T_1813_1 <= _T_584 & _T_587;
    _T_1816 <= spriteMemories_3_io_dataRead[6];
    _T_1820 <= spriteMemories_4_io_dataRead[5:0];
    _T_1822_0 <= _T_1822_1;
    if (spriteRotationReg_4) begin
      _T_1822_1 <= _T_686;
    end else begin
      _T_1822_1 <= _T_687;
    end
    _T_1825 <= spriteMemories_4_io_dataRead[6];
    _T_1829 <= spriteMemories_5_io_dataRead[5:0];
    _T_1831_0 <= _T_1831_1;
    _T_1831_1 <= _T_778 & _T_781;
    _T_1834 <= spriteMemories_5_io_dataRead[6];
    _T_1838 <= spriteMemories_6_io_dataRead[5:0];
    _T_1840_0 <= _T_1840_1;
    if (spriteRotationReg_6) begin
      _T_1840_1 <= _T_880;
    end else begin
      _T_1840_1 <= _T_881;
    end
    _T_1843 <= spriteMemories_6_io_dataRead[6];
    _T_1847 <= spriteMemories_7_io_dataRead[5:0];
    _T_1848_0 <= _T_1848_1;
    _T_1848_1 <= spriteVisibleReg_7;
    _T_1849_0 <= _T_1849_1;
    _T_1849_1 <= _T_972 & _T_975;
    _T_1852 <= spriteMemories_7_io_dataRead[6];
    _T_1856 <= spriteMemories_8_io_dataRead[5:0];
    _T_1857_0 <= _T_1857_1;
    _T_1857_1 <= spriteVisibleReg_8;
    _T_1858_0 <= _T_1858_1;
    _T_1858_1 <= _T_972 & _T_975;
    _T_1861 <= spriteMemories_8_io_dataRead[6];
    _T_1865 <= spriteMemories_9_io_dataRead[5:0];
    _T_1866_0 <= _T_1866_1;
    _T_1866_1 <= spriteVisibleReg_9;
    _T_1867_0 <= _T_1867_1;
    _T_1867_1 <= _T_972 & _T_975;
    _T_1870 <= spriteMemories_9_io_dataRead[6];
    _T_1874 <= spriteMemories_10_io_dataRead[5:0];
    _T_1875_0 <= _T_1875_1;
    _T_1875_1 <= spriteVisibleReg_10;
    _T_1876_0 <= _T_1876_1;
    _T_1876_1 <= _T_972 & _T_975;
    _T_1879 <= spriteMemories_10_io_dataRead[6];
    _T_1883 <= spriteMemories_11_io_dataRead[5:0];
    _T_1884_0 <= _T_1884_1;
    _T_1884_1 <= spriteVisibleReg_11;
    _T_1885_0 <= _T_1885_1;
    _T_1885_1 <= _T_972 & _T_975;
    _T_1888 <= spriteMemories_11_io_dataRead[6];
    _T_1892 <= spriteMemories_12_io_dataRead[5:0];
    _T_1893_0 <= _T_1893_1;
    _T_1893_1 <= spriteVisibleReg_12;
    _T_1894_0 <= _T_1894_1;
    _T_1894_1 <= _T_972 & _T_975;
    _T_1897 <= spriteMemories_12_io_dataRead[6];
    _T_1901 <= spriteMemories_13_io_dataRead[5:0];
    _T_1902_0 <= _T_1902_1;
    _T_1902_1 <= spriteVisibleReg_13;
    _T_1903_0 <= _T_1903_1;
    _T_1903_1 <= _T_972 & _T_975;
    _T_1906 <= spriteMemories_13_io_dataRead[6];
    _T_1910 <= spriteMemories_14_io_dataRead[5:0];
    _T_1911_0 <= _T_1911_1;
    _T_1911_1 <= spriteVisibleReg_14;
    _T_1912_0 <= _T_1912_1;
    _T_1912_1 <= _T_972 & _T_975;
    _T_1915 <= spriteMemories_14_io_dataRead[6];
    _T_1919 <= spriteMemories_15_io_dataRead[5:0];
    _T_1920_0 <= _T_1920_1;
    _T_1920_1 <= spriteVisibleReg_15;
    _T_1921_0 <= _T_1921_1;
    _T_1921_1 <= _T_972 & _T_975;
    _T_1924 <= spriteMemories_15_io_dataRead[6];
    pixelColorSprite <= multiHotPriortyReductionTree_io_dataOutput;
    pixelColorSpriteValid <= multiHotPriortyReductionTree_io_selectOutput;
    _T_1927_0 <= _T_1927_1;
    _T_1927_1 <= _T_1927_2;
    _T_1927_2 <= _T_17 & _T_18;
    _T_1934 <= {pixelColourVGA[5:4],pixelColourVGA[5:4]};
    _T_1935 <= {pixelColourVGA[3:2],pixelColourVGA[3:2]};
    _T_1936 <= {pixelColourVGA[1:0],pixelColourVGA[1:0]};
  end
endmodule
module Memory_51(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_52(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_53(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_54(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_55(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_56(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_57(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_58(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module SoundEngine(
  input        clock,
  input        reset,
  output       io_output_0,
  input  [3:0] io_input,
  input  [3:0] io_stop
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire  tone_0_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_0_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_0_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_1_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_1_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_1_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_2_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_2_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_2_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_3_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_3_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_3_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_4_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_4_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_4_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_5_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_5_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_5_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_6_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_6_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_6_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_7_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_7_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_7_io_dataRead; // @[SoundEngine.scala 36:23]
  reg  channel_0; // @[SoundEngine.scala 16:30]
  reg  channel_1; // @[SoundEngine.scala 16:30]
  reg  channel_2; // @[SoundEngine.scala 16:30]
  reg  channel_3; // @[SoundEngine.scala 16:30]
  reg  channel_4; // @[SoundEngine.scala 16:30]
  reg  channel_5; // @[SoundEngine.scala 16:30]
  reg  channel_6; // @[SoundEngine.scala 16:30]
  reg  channel_7; // @[SoundEngine.scala 16:30]
  reg [19:0] cntMilliSecond_0; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_1; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_2; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_3; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_4; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_5; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_6; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_7; // @[SoundEngine.scala 17:34]
  reg [19:0] slowCounter_0; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_1; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_2; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_3; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_4; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_5; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_6; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_7; // @[SoundEngine.scala 18:28]
  reg [31:0] waveCnt_0; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_1; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_2; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_3; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_4; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_5; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_6; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_7; // @[SoundEngine.scala 19:28]
  reg [8:0] toneIndex_0; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_1; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_2; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_3; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_4; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_5; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_6; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_7; // @[SoundEngine.scala 20:28]
  reg  songPlaying_0; // @[SoundEngine.scala 21:28]
  reg  songPlaying_1; // @[SoundEngine.scala 21:28]
  reg  songPlaying_2; // @[SoundEngine.scala 21:28]
  reg  songPlaying_3; // @[SoundEngine.scala 21:28]
  reg  songPlaying_4; // @[SoundEngine.scala 21:28]
  reg  songPlaying_5; // @[SoundEngine.scala 21:28]
  reg  songPlaying_6; // @[SoundEngine.scala 21:28]
  reg  songPlaying_7; // @[SoundEngine.scala 21:28]
  wire  _T_9 = io_input > 4'h0; // @[SoundEngine.scala 27:17]
  wire  _T_10 = io_input <= 4'h8; // @[SoundEngine.scala 27:35]
  wire  _T_11 = _T_9 & _T_10; // @[SoundEngine.scala 27:23]
  wire [3:0] _T_13 = io_input - 4'h1; // @[SoundEngine.scala 28:25]
  wire  _GEN_152 = 3'h0 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_8 = _GEN_152 | songPlaying_0; // @[SoundEngine.scala 28:31]
  wire  _GEN_153 = 3'h1 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_9 = _GEN_153 | songPlaying_1; // @[SoundEngine.scala 28:31]
  wire  _GEN_154 = 3'h2 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_10 = _GEN_154 | songPlaying_2; // @[SoundEngine.scala 28:31]
  wire  _GEN_155 = 3'h3 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_11 = _GEN_155 | songPlaying_3; // @[SoundEngine.scala 28:31]
  wire  _GEN_156 = 3'h4 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_12 = _GEN_156 | songPlaying_4; // @[SoundEngine.scala 28:31]
  wire  _GEN_157 = 3'h5 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_13 = _GEN_157 | songPlaying_5; // @[SoundEngine.scala 28:31]
  wire  _GEN_158 = 3'h6 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_14 = _GEN_158 | songPlaying_6; // @[SoundEngine.scala 28:31]
  wire  _GEN_159 = 3'h7 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_15 = _GEN_159 | songPlaying_7; // @[SoundEngine.scala 28:31]
  wire  _T_15 = io_stop > 4'h0; // @[SoundEngine.scala 30:16]
  wire  _T_16 = io_stop <= 4'h8; // @[SoundEngine.scala 30:33]
  wire  _T_17 = _T_15 & _T_16; // @[SoundEngine.scala 30:22]
  wire [3:0] _T_19 = io_stop - 4'h1; // @[SoundEngine.scala 31:25]
  reg [19:0] freqReg_0; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_1; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_2; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_3; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_4; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_5; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_6; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_7; // @[SoundEngine.scala 49:24]
  reg [11:0] durReg_0; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_1; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_2; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_3; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_4; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_5; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_6; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_7; // @[SoundEngine.scala 50:24]
  wire  _T_39 = ~songPlaying_0; // @[SoundEngine.scala 56:25]
  wire  _T_40 = slowCounter_0 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_42 = cntMilliSecond_0 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_44 = slowCounter_0 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_45 = freqReg_0 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_47 = waveCnt_0 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_160 = {{12'd0}, freqReg_0}; // @[SoundEngine.scala 81:23]
  wire  _T_48 = waveCnt_0 >= _GEN_160; // @[SoundEngine.scala 81:23]
  wire  _T_49 = ~channel_0; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_161 = {{8'd0}, durReg_0}; // @[SoundEngine.scala 88:28]
  wire  _T_50 = cntMilliSecond_0 >= _GEN_161; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_52 = toneIndex_0 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_53 = durReg_0 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_54 = ~songPlaying_1; // @[SoundEngine.scala 56:25]
  wire  _T_55 = slowCounter_1 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_57 = cntMilliSecond_1 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_59 = slowCounter_1 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_60 = freqReg_1 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_62 = waveCnt_1 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_162 = {{12'd0}, freqReg_1}; // @[SoundEngine.scala 81:23]
  wire  _T_63 = waveCnt_1 >= _GEN_162; // @[SoundEngine.scala 81:23]
  wire  _T_64 = ~channel_1; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_163 = {{8'd0}, durReg_1}; // @[SoundEngine.scala 88:28]
  wire  _T_65 = cntMilliSecond_1 >= _GEN_163; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_67 = toneIndex_1 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_68 = durReg_1 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_69 = ~songPlaying_2; // @[SoundEngine.scala 56:25]
  wire  _T_70 = slowCounter_2 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_72 = cntMilliSecond_2 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_74 = slowCounter_2 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_75 = freqReg_2 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_77 = waveCnt_2 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_164 = {{12'd0}, freqReg_2}; // @[SoundEngine.scala 81:23]
  wire  _T_78 = waveCnt_2 >= _GEN_164; // @[SoundEngine.scala 81:23]
  wire  _T_79 = ~channel_2; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_165 = {{8'd0}, durReg_2}; // @[SoundEngine.scala 88:28]
  wire  _T_80 = cntMilliSecond_2 >= _GEN_165; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_82 = toneIndex_2 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_83 = durReg_2 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_84 = ~songPlaying_3; // @[SoundEngine.scala 56:25]
  wire  _T_85 = slowCounter_3 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_87 = cntMilliSecond_3 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_89 = slowCounter_3 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_90 = freqReg_3 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_92 = waveCnt_3 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_166 = {{12'd0}, freqReg_3}; // @[SoundEngine.scala 81:23]
  wire  _T_93 = waveCnt_3 >= _GEN_166; // @[SoundEngine.scala 81:23]
  wire  _T_94 = ~channel_3; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_167 = {{8'd0}, durReg_3}; // @[SoundEngine.scala 88:28]
  wire  _T_95 = cntMilliSecond_3 >= _GEN_167; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_97 = toneIndex_3 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_98 = durReg_3 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_99 = ~songPlaying_4; // @[SoundEngine.scala 56:25]
  wire  _T_100 = slowCounter_4 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_102 = cntMilliSecond_4 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_104 = slowCounter_4 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_105 = freqReg_4 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_107 = waveCnt_4 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_168 = {{12'd0}, freqReg_4}; // @[SoundEngine.scala 81:23]
  wire  _T_108 = waveCnt_4 >= _GEN_168; // @[SoundEngine.scala 81:23]
  wire  _T_109 = ~channel_4; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_169 = {{8'd0}, durReg_4}; // @[SoundEngine.scala 88:28]
  wire  _T_110 = cntMilliSecond_4 >= _GEN_169; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_112 = toneIndex_4 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_113 = durReg_4 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_114 = ~songPlaying_5; // @[SoundEngine.scala 56:25]
  wire  _T_115 = slowCounter_5 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_117 = cntMilliSecond_5 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_119 = slowCounter_5 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_120 = freqReg_5 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_122 = waveCnt_5 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_170 = {{12'd0}, freqReg_5}; // @[SoundEngine.scala 81:23]
  wire  _T_123 = waveCnt_5 >= _GEN_170; // @[SoundEngine.scala 81:23]
  wire  _T_124 = ~channel_5; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_171 = {{8'd0}, durReg_5}; // @[SoundEngine.scala 88:28]
  wire  _T_125 = cntMilliSecond_5 >= _GEN_171; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_127 = toneIndex_5 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_128 = durReg_5 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_129 = ~songPlaying_6; // @[SoundEngine.scala 56:25]
  wire  _T_130 = slowCounter_6 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_132 = cntMilliSecond_6 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_134 = slowCounter_6 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_135 = freqReg_6 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_137 = waveCnt_6 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_172 = {{12'd0}, freqReg_6}; // @[SoundEngine.scala 81:23]
  wire  _T_138 = waveCnt_6 >= _GEN_172; // @[SoundEngine.scala 81:23]
  wire  _T_139 = ~channel_6; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_173 = {{8'd0}, durReg_6}; // @[SoundEngine.scala 88:28]
  wire  _T_140 = cntMilliSecond_6 >= _GEN_173; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_142 = toneIndex_6 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_143 = durReg_6 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_144 = ~songPlaying_7; // @[SoundEngine.scala 56:25]
  wire  _T_145 = slowCounter_7 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_147 = cntMilliSecond_7 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_149 = slowCounter_7 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_150 = freqReg_7 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_152 = waveCnt_7 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_174 = {{12'd0}, freqReg_7}; // @[SoundEngine.scala 81:23]
  wire  _T_153 = waveCnt_7 >= _GEN_174; // @[SoundEngine.scala 81:23]
  wire  _T_154 = ~channel_7; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_175 = {{8'd0}, durReg_7}; // @[SoundEngine.scala 88:28]
  wire  _T_155 = cntMilliSecond_7 >= _GEN_175; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_157 = toneIndex_7 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_158 = durReg_7 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_159 = channel_0 | channel_1; // @[SoundEngine.scala 98:35]
  wire  _T_160 = _T_159 | channel_2; // @[SoundEngine.scala 98:35]
  wire  _T_161 = _T_160 | channel_3; // @[SoundEngine.scala 98:35]
  wire  _T_162 = _T_161 | channel_4; // @[SoundEngine.scala 98:35]
  wire  _T_163 = _T_162 | channel_5; // @[SoundEngine.scala 98:35]
  wire  _T_164 = _T_163 | channel_6; // @[SoundEngine.scala 98:35]
  Memory_51 tone_0 ( // @[SoundEngine.scala 36:23]
    .clock(tone_0_clock),
    .io_address(tone_0_io_address),
    .io_dataRead(tone_0_io_dataRead)
  );
  Memory_52 tone_1 ( // @[SoundEngine.scala 36:23]
    .clock(tone_1_clock),
    .io_address(tone_1_io_address),
    .io_dataRead(tone_1_io_dataRead)
  );
  Memory_53 tone_2 ( // @[SoundEngine.scala 36:23]
    .clock(tone_2_clock),
    .io_address(tone_2_io_address),
    .io_dataRead(tone_2_io_dataRead)
  );
  Memory_54 tone_3 ( // @[SoundEngine.scala 36:23]
    .clock(tone_3_clock),
    .io_address(tone_3_io_address),
    .io_dataRead(tone_3_io_dataRead)
  );
  Memory_55 tone_4 ( // @[SoundEngine.scala 36:23]
    .clock(tone_4_clock),
    .io_address(tone_4_io_address),
    .io_dataRead(tone_4_io_dataRead)
  );
  Memory_56 tone_5 ( // @[SoundEngine.scala 36:23]
    .clock(tone_5_clock),
    .io_address(tone_5_io_address),
    .io_dataRead(tone_5_io_dataRead)
  );
  Memory_57 tone_6 ( // @[SoundEngine.scala 36:23]
    .clock(tone_6_clock),
    .io_address(tone_6_io_address),
    .io_dataRead(tone_6_io_dataRead)
  );
  Memory_58 tone_7 ( // @[SoundEngine.scala 36:23]
    .clock(tone_7_clock),
    .io_address(tone_7_io_address),
    .io_dataRead(tone_7_io_dataRead)
  );
  assign io_output_0 = _T_164 | channel_7; // @[SoundEngine.scala 98:16]
  assign tone_0_clock = clock;
  assign tone_0_io_address = toneIndex_0; // @[SoundEngine.scala 45:24]
  assign tone_1_clock = clock;
  assign tone_1_io_address = toneIndex_1; // @[SoundEngine.scala 45:24]
  assign tone_2_clock = clock;
  assign tone_2_io_address = toneIndex_2; // @[SoundEngine.scala 45:24]
  assign tone_3_clock = clock;
  assign tone_3_io_address = toneIndex_3; // @[SoundEngine.scala 45:24]
  assign tone_4_clock = clock;
  assign tone_4_io_address = toneIndex_4; // @[SoundEngine.scala 45:24]
  assign tone_5_clock = clock;
  assign tone_5_io_address = toneIndex_5; // @[SoundEngine.scala 45:24]
  assign tone_6_clock = clock;
  assign tone_6_io_address = toneIndex_6; // @[SoundEngine.scala 45:24]
  assign tone_7_clock = clock;
  assign tone_7_io_address = toneIndex_7; // @[SoundEngine.scala 45:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  channel_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  channel_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  channel_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  channel_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  channel_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  channel_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  channel_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  channel_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cntMilliSecond_0 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  cntMilliSecond_1 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  cntMilliSecond_2 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  cntMilliSecond_3 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  cntMilliSecond_4 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  cntMilliSecond_5 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  cntMilliSecond_6 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  cntMilliSecond_7 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  slowCounter_0 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  slowCounter_1 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  slowCounter_2 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  slowCounter_3 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  slowCounter_4 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  slowCounter_5 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  slowCounter_6 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  slowCounter_7 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  waveCnt_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  waveCnt_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  waveCnt_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  waveCnt_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  waveCnt_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  waveCnt_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  waveCnt_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  waveCnt_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  toneIndex_0 = _RAND_32[8:0];
  _RAND_33 = {1{`RANDOM}};
  toneIndex_1 = _RAND_33[8:0];
  _RAND_34 = {1{`RANDOM}};
  toneIndex_2 = _RAND_34[8:0];
  _RAND_35 = {1{`RANDOM}};
  toneIndex_3 = _RAND_35[8:0];
  _RAND_36 = {1{`RANDOM}};
  toneIndex_4 = _RAND_36[8:0];
  _RAND_37 = {1{`RANDOM}};
  toneIndex_5 = _RAND_37[8:0];
  _RAND_38 = {1{`RANDOM}};
  toneIndex_6 = _RAND_38[8:0];
  _RAND_39 = {1{`RANDOM}};
  toneIndex_7 = _RAND_39[8:0];
  _RAND_40 = {1{`RANDOM}};
  songPlaying_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  songPlaying_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  songPlaying_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  songPlaying_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  songPlaying_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  songPlaying_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  songPlaying_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  songPlaying_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  freqReg_0 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  freqReg_1 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  freqReg_2 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  freqReg_3 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  freqReg_4 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  freqReg_5 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  freqReg_6 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  freqReg_7 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  durReg_0 = _RAND_56[11:0];
  _RAND_57 = {1{`RANDOM}};
  durReg_1 = _RAND_57[11:0];
  _RAND_58 = {1{`RANDOM}};
  durReg_2 = _RAND_58[11:0];
  _RAND_59 = {1{`RANDOM}};
  durReg_3 = _RAND_59[11:0];
  _RAND_60 = {1{`RANDOM}};
  durReg_4 = _RAND_60[11:0];
  _RAND_61 = {1{`RANDOM}};
  durReg_5 = _RAND_61[11:0];
  _RAND_62 = {1{`RANDOM}};
  durReg_6 = _RAND_62[11:0];
  _RAND_63 = {1{`RANDOM}};
  durReg_7 = _RAND_63[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      channel_0 <= 1'h0;
    end else if (_T_45) begin
      channel_0 <= 1'h0;
    end else if (_T_48) begin
      channel_0 <= _T_49;
    end else if (_T_39) begin
      channel_0 <= 1'h0;
    end
    if (reset) begin
      channel_1 <= 1'h0;
    end else if (_T_60) begin
      channel_1 <= 1'h0;
    end else if (_T_63) begin
      channel_1 <= _T_64;
    end else if (_T_54) begin
      channel_1 <= 1'h0;
    end
    if (reset) begin
      channel_2 <= 1'h0;
    end else if (_T_75) begin
      channel_2 <= 1'h0;
    end else if (_T_78) begin
      channel_2 <= _T_79;
    end else if (_T_69) begin
      channel_2 <= 1'h0;
    end
    if (reset) begin
      channel_3 <= 1'h0;
    end else if (_T_90) begin
      channel_3 <= 1'h0;
    end else if (_T_93) begin
      channel_3 <= _T_94;
    end else if (_T_84) begin
      channel_3 <= 1'h0;
    end
    if (reset) begin
      channel_4 <= 1'h0;
    end else if (_T_105) begin
      channel_4 <= 1'h0;
    end else if (_T_108) begin
      channel_4 <= _T_109;
    end else if (_T_99) begin
      channel_4 <= 1'h0;
    end
    if (reset) begin
      channel_5 <= 1'h0;
    end else if (_T_120) begin
      channel_5 <= 1'h0;
    end else if (_T_123) begin
      channel_5 <= _T_124;
    end else if (_T_114) begin
      channel_5 <= 1'h0;
    end
    if (reset) begin
      channel_6 <= 1'h0;
    end else if (_T_135) begin
      channel_6 <= 1'h0;
    end else if (_T_138) begin
      channel_6 <= _T_139;
    end else if (_T_129) begin
      channel_6 <= 1'h0;
    end
    if (reset) begin
      channel_7 <= 1'h0;
    end else if (_T_150) begin
      channel_7 <= 1'h0;
    end else if (_T_153) begin
      channel_7 <= _T_154;
    end else if (_T_144) begin
      channel_7 <= 1'h0;
    end
    if (reset) begin
      cntMilliSecond_0 <= 20'h0;
    end else if (_T_50) begin
      cntMilliSecond_0 <= 20'h0;
    end else if (_T_40) begin
      cntMilliSecond_0 <= _T_42;
    end else if (_T_39) begin
      cntMilliSecond_0 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_1 <= 20'h0;
    end else if (_T_65) begin
      cntMilliSecond_1 <= 20'h0;
    end else if (_T_55) begin
      cntMilliSecond_1 <= _T_57;
    end else if (_T_54) begin
      cntMilliSecond_1 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_2 <= 20'h0;
    end else if (_T_80) begin
      cntMilliSecond_2 <= 20'h0;
    end else if (_T_70) begin
      cntMilliSecond_2 <= _T_72;
    end else if (_T_69) begin
      cntMilliSecond_2 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_3 <= 20'h0;
    end else if (_T_95) begin
      cntMilliSecond_3 <= 20'h0;
    end else if (_T_85) begin
      cntMilliSecond_3 <= _T_87;
    end else if (_T_84) begin
      cntMilliSecond_3 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_4 <= 20'h0;
    end else if (_T_110) begin
      cntMilliSecond_4 <= 20'h0;
    end else if (_T_100) begin
      cntMilliSecond_4 <= _T_102;
    end else if (_T_99) begin
      cntMilliSecond_4 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_5 <= 20'h0;
    end else if (_T_125) begin
      cntMilliSecond_5 <= 20'h0;
    end else if (_T_115) begin
      cntMilliSecond_5 <= _T_117;
    end else if (_T_114) begin
      cntMilliSecond_5 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_6 <= 20'h0;
    end else if (_T_140) begin
      cntMilliSecond_6 <= 20'h0;
    end else if (_T_130) begin
      cntMilliSecond_6 <= _T_132;
    end else if (_T_129) begin
      cntMilliSecond_6 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_7 <= 20'h0;
    end else if (_T_155) begin
      cntMilliSecond_7 <= 20'h0;
    end else if (_T_145) begin
      cntMilliSecond_7 <= _T_147;
    end else if (_T_144) begin
      cntMilliSecond_7 <= 20'h0;
    end
    if (reset) begin
      slowCounter_0 <= 20'h0;
    end else if (_T_40) begin
      slowCounter_0 <= 20'h0;
    end else begin
      slowCounter_0 <= _T_44;
    end
    if (reset) begin
      slowCounter_1 <= 20'h0;
    end else if (_T_55) begin
      slowCounter_1 <= 20'h0;
    end else begin
      slowCounter_1 <= _T_59;
    end
    if (reset) begin
      slowCounter_2 <= 20'h0;
    end else if (_T_70) begin
      slowCounter_2 <= 20'h0;
    end else begin
      slowCounter_2 <= _T_74;
    end
    if (reset) begin
      slowCounter_3 <= 20'h0;
    end else if (_T_85) begin
      slowCounter_3 <= 20'h0;
    end else begin
      slowCounter_3 <= _T_89;
    end
    if (reset) begin
      slowCounter_4 <= 20'h0;
    end else if (_T_100) begin
      slowCounter_4 <= 20'h0;
    end else begin
      slowCounter_4 <= _T_104;
    end
    if (reset) begin
      slowCounter_5 <= 20'h0;
    end else if (_T_115) begin
      slowCounter_5 <= 20'h0;
    end else begin
      slowCounter_5 <= _T_119;
    end
    if (reset) begin
      slowCounter_6 <= 20'h0;
    end else if (_T_130) begin
      slowCounter_6 <= 20'h0;
    end else begin
      slowCounter_6 <= _T_134;
    end
    if (reset) begin
      slowCounter_7 <= 20'h0;
    end else if (_T_145) begin
      slowCounter_7 <= 20'h0;
    end else begin
      slowCounter_7 <= _T_149;
    end
    if (reset) begin
      waveCnt_0 <= 32'h0;
    end else if (_T_45) begin
      waveCnt_0 <= 32'h0;
    end else if (_T_48) begin
      waveCnt_0 <= 32'h0;
    end else begin
      waveCnt_0 <= _T_47;
    end
    if (reset) begin
      waveCnt_1 <= 32'h0;
    end else if (_T_60) begin
      waveCnt_1 <= 32'h0;
    end else if (_T_63) begin
      waveCnt_1 <= 32'h0;
    end else begin
      waveCnt_1 <= _T_62;
    end
    if (reset) begin
      waveCnt_2 <= 32'h0;
    end else if (_T_75) begin
      waveCnt_2 <= 32'h0;
    end else if (_T_78) begin
      waveCnt_2 <= 32'h0;
    end else begin
      waveCnt_2 <= _T_77;
    end
    if (reset) begin
      waveCnt_3 <= 32'h0;
    end else if (_T_90) begin
      waveCnt_3 <= 32'h0;
    end else if (_T_93) begin
      waveCnt_3 <= 32'h0;
    end else begin
      waveCnt_3 <= _T_92;
    end
    if (reset) begin
      waveCnt_4 <= 32'h0;
    end else if (_T_105) begin
      waveCnt_4 <= 32'h0;
    end else if (_T_108) begin
      waveCnt_4 <= 32'h0;
    end else begin
      waveCnt_4 <= _T_107;
    end
    if (reset) begin
      waveCnt_5 <= 32'h0;
    end else if (_T_120) begin
      waveCnt_5 <= 32'h0;
    end else if (_T_123) begin
      waveCnt_5 <= 32'h0;
    end else begin
      waveCnt_5 <= _T_122;
    end
    if (reset) begin
      waveCnt_6 <= 32'h0;
    end else if (_T_135) begin
      waveCnt_6 <= 32'h0;
    end else if (_T_138) begin
      waveCnt_6 <= 32'h0;
    end else begin
      waveCnt_6 <= _T_137;
    end
    if (reset) begin
      waveCnt_7 <= 32'h0;
    end else if (_T_150) begin
      waveCnt_7 <= 32'h0;
    end else if (_T_153) begin
      waveCnt_7 <= 32'h0;
    end else begin
      waveCnt_7 <= _T_152;
    end
    if (reset) begin
      toneIndex_0 <= 9'h0;
    end else if (_T_50) begin
      toneIndex_0 <= _T_52;
    end else if (_T_39) begin
      toneIndex_0 <= 9'h0;
    end
    if (reset) begin
      toneIndex_1 <= 9'h0;
    end else if (_T_65) begin
      toneIndex_1 <= _T_67;
    end else if (_T_54) begin
      toneIndex_1 <= 9'h0;
    end
    if (reset) begin
      toneIndex_2 <= 9'h0;
    end else if (_T_80) begin
      toneIndex_2 <= _T_82;
    end else if (_T_69) begin
      toneIndex_2 <= 9'h0;
    end
    if (reset) begin
      toneIndex_3 <= 9'h0;
    end else if (_T_95) begin
      toneIndex_3 <= _T_97;
    end else if (_T_84) begin
      toneIndex_3 <= 9'h0;
    end
    if (reset) begin
      toneIndex_4 <= 9'h0;
    end else if (_T_110) begin
      toneIndex_4 <= _T_112;
    end else if (_T_99) begin
      toneIndex_4 <= 9'h0;
    end
    if (reset) begin
      toneIndex_5 <= 9'h0;
    end else if (_T_125) begin
      toneIndex_5 <= _T_127;
    end else if (_T_114) begin
      toneIndex_5 <= 9'h0;
    end
    if (reset) begin
      toneIndex_6 <= 9'h0;
    end else if (_T_140) begin
      toneIndex_6 <= _T_142;
    end else if (_T_129) begin
      toneIndex_6 <= 9'h0;
    end
    if (reset) begin
      toneIndex_7 <= 9'h0;
    end else if (_T_155) begin
      toneIndex_7 <= _T_157;
    end else if (_T_144) begin
      toneIndex_7 <= 9'h0;
    end
    if (reset) begin
      songPlaying_0 <= 1'h0;
    end else if (_T_53) begin
      songPlaying_0 <= 1'h0;
    end else if (_T_17) begin
      if (3'h0 == _T_19[2:0]) begin
        songPlaying_0 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_0 <= _GEN_8;
      end
    end else if (_T_11) begin
      songPlaying_0 <= _GEN_8;
    end
    if (reset) begin
      songPlaying_1 <= 1'h0;
    end else if (_T_68) begin
      songPlaying_1 <= 1'h0;
    end else if (_T_17) begin
      if (3'h1 == _T_19[2:0]) begin
        songPlaying_1 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_1 <= _GEN_9;
      end
    end else if (_T_11) begin
      songPlaying_1 <= _GEN_9;
    end
    if (reset) begin
      songPlaying_2 <= 1'h0;
    end else if (_T_83) begin
      songPlaying_2 <= 1'h0;
    end else if (_T_17) begin
      if (3'h2 == _T_19[2:0]) begin
        songPlaying_2 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_2 <= _GEN_10;
      end
    end else if (_T_11) begin
      songPlaying_2 <= _GEN_10;
    end
    if (reset) begin
      songPlaying_3 <= 1'h0;
    end else if (_T_98) begin
      songPlaying_3 <= 1'h0;
    end else if (_T_17) begin
      if (3'h3 == _T_19[2:0]) begin
        songPlaying_3 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_3 <= _GEN_11;
      end
    end else if (_T_11) begin
      songPlaying_3 <= _GEN_11;
    end
    if (reset) begin
      songPlaying_4 <= 1'h0;
    end else if (_T_113) begin
      songPlaying_4 <= 1'h0;
    end else if (_T_17) begin
      if (3'h4 == _T_19[2:0]) begin
        songPlaying_4 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_4 <= _GEN_12;
      end
    end else if (_T_11) begin
      songPlaying_4 <= _GEN_12;
    end
    if (reset) begin
      songPlaying_5 <= 1'h0;
    end else if (_T_128) begin
      songPlaying_5 <= 1'h0;
    end else if (_T_17) begin
      if (3'h5 == _T_19[2:0]) begin
        songPlaying_5 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_5 <= _GEN_13;
      end
    end else if (_T_11) begin
      songPlaying_5 <= _GEN_13;
    end
    if (reset) begin
      songPlaying_6 <= 1'h0;
    end else if (_T_143) begin
      songPlaying_6 <= 1'h0;
    end else if (_T_17) begin
      if (3'h6 == _T_19[2:0]) begin
        songPlaying_6 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_6 <= _GEN_14;
      end
    end else if (_T_11) begin
      songPlaying_6 <= _GEN_14;
    end
    if (reset) begin
      songPlaying_7 <= 1'h0;
    end else if (_T_158) begin
      songPlaying_7 <= 1'h0;
    end else if (_T_17) begin
      if (3'h7 == _T_19[2:0]) begin
        songPlaying_7 <= 1'h0;
      end else if (_T_11) begin
        songPlaying_7 <= _GEN_15;
      end
    end else if (_T_11) begin
      songPlaying_7 <= _GEN_15;
    end
    freqReg_0 <= tone_0_io_dataRead[31:12];
    freqReg_1 <= tone_1_io_dataRead[31:12];
    freqReg_2 <= tone_2_io_dataRead[31:12];
    freqReg_3 <= tone_3_io_dataRead[31:12];
    freqReg_4 <= tone_4_io_dataRead[31:12];
    freqReg_5 <= tone_5_io_dataRead[31:12];
    freqReg_6 <= tone_6_io_dataRead[31:12];
    freqReg_7 <= tone_7_io_dataRead[31:12];
    durReg_0 <= tone_0_io_dataRead[11:0];
    durReg_1 <= tone_1_io_dataRead[11:0];
    durReg_2 <= tone_2_io_dataRead[11:0];
    durReg_3 <= tone_3_io_dataRead[11:0];
    durReg_4 <= tone_4_io_dataRead[11:0];
    durReg_5 <= tone_5_io_dataRead[11:0];
    durReg_6 <= tone_6_io_dataRead[11:0];
    durReg_7 <= tone_7_io_dataRead[11:0];
  end
endmodule
module GameLogicTask3(
  input         clock,
  input         reset,
  input         io_btnC,
  input         io_btnU,
  input         io_btnL,
  input         io_btnR,
  input         io_btnD,
  output [3:0]  io_songInput,
  output [3:0]  io_songStop,
  output [10:0] io_spriteXPosition_0,
  output [9:0]  io_spriteYPosition_0,
  output        io_spriteFlipHorizontal_0,
  input         io_newFrame,
  output        io_frameUpdateDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[GameLogicTask3.scala 109:25]
  reg [10:0] sprite0XReg; // @[GameLogicTask3.scala 112:28]
  reg [9:0] sprite0YReg; // @[GameLogicTask3.scala 113:28]
  reg  sprite0FlipHorizontalReg; // @[GameLogicTask3.scala 116:41]
  wire  _T = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = $signed(sprite0YReg) < 10'sh1a8; // @[GameLogicTask3.scala 192:26]
  wire [9:0] _T_5 = $signed(sprite0YReg) + 10'sh2; // @[GameLogicTask3.scala 193:38]
  wire  _GEN_2 = _T_2 ? 1'h0 : sprite0FlipHorizontalReg; // @[GameLogicTask3.scala 192:47]
  wire [1:0] _GEN_3 = _T_2 ? 2'h3 : 2'h0; // @[GameLogicTask3.scala 192:47]
  wire  _T_6 = $signed(sprite0YReg) > 10'sh60; // @[GameLogicTask3.scala 199:26]
  wire [9:0] _T_9 = $signed(sprite0YReg) - 10'sh2; // @[GameLogicTask3.scala 200:38]
  wire  _GEN_5 = _T_6 | sprite0FlipHorizontalReg; // @[GameLogicTask3.scala 199:36]
  wire [1:0] _GEN_6 = _T_6 ? 2'h2 : 2'h0; // @[GameLogicTask3.scala 199:36]
  wire  _GEN_8 = io_btnU ? _GEN_5 : sprite0FlipHorizontalReg; // @[GameLogicTask3.scala 198:27]
  wire [1:0] _GEN_9 = io_btnU ? _GEN_6 : 2'h0; // @[GameLogicTask3.scala 198:27]
  wire  _GEN_11 = io_btnD ? _GEN_2 : _GEN_8; // @[GameLogicTask3.scala 191:20]
  wire [1:0] _GEN_12 = io_btnD ? _GEN_3 : _GEN_9; // @[GameLogicTask3.scala 191:20]
  wire [1:0] _GEN_13 = io_btnC ? 2'h1 : _GEN_12; // @[GameLogicTask3.scala 208:20]
  wire  _T_10 = $signed(sprite0XReg) < 11'sh240; // @[GameLogicTask3.scala 212:26]
  wire [10:0] _T_13 = $signed(sprite0XReg) + 11'sh2; // @[GameLogicTask3.scala 213:38]
  wire [2:0] _GEN_16 = _T_10 ? 3'h4 : {{1'd0}, _GEN_13}; // @[GameLogicTask3.scala 212:47]
  wire  _T_14 = $signed(sprite0XReg) > 11'sh20; // @[GameLogicTask3.scala 219:26]
  wire [10:0] _T_17 = $signed(sprite0XReg) - 11'sh2; // @[GameLogicTask3.scala 220:38]
  wire  _GEN_18 = _T_14 | _GEN_11; // @[GameLogicTask3.scala 219:34]
  wire [1:0] _GEN_19 = _T_14 ? 2'h2 : 2'h0; // @[GameLogicTask3.scala 219:34]
  wire [1:0] _GEN_22 = io_btnL ? _GEN_19 : 2'h0; // @[GameLogicTask3.scala 218:27]
  wire [2:0] _GEN_25 = io_btnR ? _GEN_16 : {{1'd0}, _GEN_13}; // @[GameLogicTask3.scala 211:21]
  wire [1:0] _GEN_26 = io_btnR ? 2'h0 : _GEN_22; // @[GameLogicTask3.scala 211:21]
  wire  _T_18 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_31 = _T_1 ? _GEN_25 : 3'h0; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_33 = _T_1 ? _GEN_26 : 2'h0; // @[Conditional.scala 39:67]
  wire  _GEN_35 = _T_1 ? 1'h0 : _T_18; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_39 = _T ? 3'h0 : _GEN_31; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_41 = _T ? 2'h0 : _GEN_33; // @[Conditional.scala 40:58]
  assign io_songInput = {{1'd0}, _GEN_39}; // @[GameLogicTask3.scala 88:14 GameLogicTask3.scala 195:23 GameLogicTask3.scala 202:23 GameLogicTask3.scala 209:21 GameLogicTask3.scala 215:23]
  assign io_songStop = {{2'd0}, _GEN_41}; // @[GameLogicTask3.scala 89:14 GameLogicTask3.scala 222:22]
  assign io_spriteXPosition_0 = sprite0XReg; // @[GameLogicTask3.scala 79:22 GameLogicTask3.scala 173:25]
  assign io_spriteYPosition_0 = sprite0YReg; // @[GameLogicTask3.scala 80:22 GameLogicTask3.scala 174:25]
  assign io_spriteFlipHorizontal_0 = sprite0FlipHorizontalReg; // @[GameLogicTask3.scala 82:27 GameLogicTask3.scala 175:30]
  assign io_frameUpdateDone = _T ? 1'h0 : _GEN_35; // @[GameLogicTask3.scala 104:22 GameLogicTask3.scala 244:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  sprite0XReg = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  sprite0YReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  sprite0FlipHorizontalReg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T) begin
      if (io_newFrame) begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      stateReg <= 2'h2;
    end else if (_T_18) begin
      stateReg <= 2'h0;
    end
    if (reset) begin
      sprite0XReg <= 11'sh20;
    end else if (!(_T)) begin
      if (_T_1) begin
        if (io_btnR) begin
          if (_T_10) begin
            sprite0XReg <= _T_13;
          end
        end else if (io_btnL) begin
          if (_T_14) begin
            sprite0XReg <= _T_17;
          end
        end
      end
    end
    if (reset) begin
      sprite0YReg <= 10'sh148;
    end else if (!(_T)) begin
      if (_T_1) begin
        if (io_btnD) begin
          if (_T_2) begin
            sprite0YReg <= _T_5;
          end
        end else if (io_btnU) begin
          if (_T_6) begin
            sprite0YReg <= _T_9;
          end
        end
      end
    end
    if (reset) begin
      sprite0FlipHorizontalReg <= 1'h0;
    end else if (!(_T)) begin
      if (_T_1) begin
        if (io_btnR) begin
          if (_T_10) begin
            sprite0FlipHorizontalReg <= 1'h0;
          end else if (io_btnD) begin
            if (_T_2) begin
              sprite0FlipHorizontalReg <= 1'h0;
            end
          end else if (io_btnU) begin
            sprite0FlipHorizontalReg <= _GEN_5;
          end
        end else if (io_btnL) begin
          sprite0FlipHorizontalReg <= _GEN_18;
        end else if (io_btnD) begin
          if (_T_2) begin
            sprite0FlipHorizontalReg <= 1'h0;
          end
        end else if (io_btnU) begin
          sprite0FlipHorizontalReg <= _GEN_5;
        end
      end
    end
  end
endmodule
module GameTop(
  input        clock,
  input        reset,
  input        io_btnC,
  input        io_btnU,
  input        io_btnL,
  input        io_btnR,
  input        io_btnD,
  output [3:0] io_vgaRed,
  output [3:0] io_vgaBlue,
  output [3:0] io_vgaGreen,
  output       io_Hsync,
  output       io_Vsync,
  output       io_soundOutput_0,
  output       io_missingFrameError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  graphicEngineVGA_clock; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_reset; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_0; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_0; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipHorizontal_0; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_newFrame; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_frameUpdateDone; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_missingFrameError; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaRed; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaBlue; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaGreen; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Hsync; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Vsync; // @[GameTop.scala 46:32]
  wire  soundEngine_clock; // @[GameTop.scala 48:27]
  wire  soundEngine_reset; // @[GameTop.scala 48:27]
  wire  soundEngine_io_output_0; // @[GameTop.scala 48:27]
  wire [3:0] soundEngine_io_input; // @[GameTop.scala 48:27]
  wire [3:0] soundEngine_io_stop; // @[GameTop.scala 48:27]
  wire  gameLogic_clock; // @[GameTop.scala 56:25]
  wire  gameLogic_reset; // @[GameTop.scala 56:25]
  wire  gameLogic_io_btnC; // @[GameTop.scala 56:25]
  wire  gameLogic_io_btnU; // @[GameTop.scala 56:25]
  wire  gameLogic_io_btnL; // @[GameTop.scala 56:25]
  wire  gameLogic_io_btnR; // @[GameTop.scala 56:25]
  wire  gameLogic_io_btnD; // @[GameTop.scala 56:25]
  wire [3:0] gameLogic_io_songInput; // @[GameTop.scala 56:25]
  wire [3:0] gameLogic_io_songStop; // @[GameTop.scala 56:25]
  wire [10:0] gameLogic_io_spriteXPosition_0; // @[GameTop.scala 56:25]
  wire [9:0] gameLogic_io_spriteYPosition_0; // @[GameTop.scala 56:25]
  wire  gameLogic_io_spriteFlipHorizontal_0; // @[GameTop.scala 56:25]
  wire  gameLogic_io_newFrame; // @[GameTop.scala 56:25]
  wire  gameLogic_io_frameUpdateDone; // @[GameTop.scala 56:25]
  reg [20:0] debounceCounter; // @[GameTop.scala 67:32]
  wire  debounceSampleEn = debounceCounter == 21'h1e847f; // @[GameTop.scala 69:24]
  wire [20:0] _T_2 = debounceCounter + 21'h1; // @[GameTop.scala 73:40]
  reg [21:0] resetReleaseCounter; // @[GameTop.scala 80:36]
  wire  _T_3 = resetReleaseCounter == 22'h3d08ff; // @[GameTop.scala 82:28]
  wire [21:0] _T_5 = resetReleaseCounter + 22'h1; // @[GameTop.scala 86:48]
  reg  _T_7_0; // @[GameUtilities.scala 39:28]
  reg  _T_7_1; // @[GameUtilities.scala 39:28]
  reg  _T_7_2; // @[GameUtilities.scala 39:28]
  reg  btnCState; // @[Reg.scala 27:20]
  reg  _T_9_0; // @[GameUtilities.scala 39:28]
  reg  _T_9_1; // @[GameUtilities.scala 39:28]
  reg  _T_9_2; // @[GameUtilities.scala 39:28]
  reg  btnUState; // @[Reg.scala 27:20]
  reg  _T_11_0; // @[GameUtilities.scala 39:28]
  reg  _T_11_1; // @[GameUtilities.scala 39:28]
  reg  _T_11_2; // @[GameUtilities.scala 39:28]
  reg  btnLState; // @[Reg.scala 27:20]
  reg  _T_13_0; // @[GameUtilities.scala 39:28]
  reg  _T_13_1; // @[GameUtilities.scala 39:28]
  reg  _T_13_2; // @[GameUtilities.scala 39:28]
  reg  btnRState; // @[Reg.scala 27:20]
  reg  _T_15_0; // @[GameUtilities.scala 39:28]
  reg  _T_15_1; // @[GameUtilities.scala 39:28]
  reg  _T_15_2; // @[GameUtilities.scala 39:28]
  reg  btnDState; // @[Reg.scala 27:20]
  GraphicEngineVGA graphicEngineVGA ( // @[GameTop.scala 46:32]
    .clock(graphicEngineVGA_clock),
    .reset(graphicEngineVGA_reset),
    .io_spriteXPosition_0(graphicEngineVGA_io_spriteXPosition_0),
    .io_spriteYPosition_0(graphicEngineVGA_io_spriteYPosition_0),
    .io_spriteFlipHorizontal_0(graphicEngineVGA_io_spriteFlipHorizontal_0),
    .io_newFrame(graphicEngineVGA_io_newFrame),
    .io_frameUpdateDone(graphicEngineVGA_io_frameUpdateDone),
    .io_missingFrameError(graphicEngineVGA_io_missingFrameError),
    .io_vgaRed(graphicEngineVGA_io_vgaRed),
    .io_vgaBlue(graphicEngineVGA_io_vgaBlue),
    .io_vgaGreen(graphicEngineVGA_io_vgaGreen),
    .io_Hsync(graphicEngineVGA_io_Hsync),
    .io_Vsync(graphicEngineVGA_io_Vsync)
  );
  SoundEngine soundEngine ( // @[GameTop.scala 48:27]
    .clock(soundEngine_clock),
    .reset(soundEngine_reset),
    .io_output_0(soundEngine_io_output_0),
    .io_input(soundEngine_io_input),
    .io_stop(soundEngine_io_stop)
  );
  GameLogicTask3 gameLogic ( // @[GameTop.scala 56:25]
    .clock(gameLogic_clock),
    .reset(gameLogic_reset),
    .io_btnC(gameLogic_io_btnC),
    .io_btnU(gameLogic_io_btnU),
    .io_btnL(gameLogic_io_btnL),
    .io_btnR(gameLogic_io_btnR),
    .io_btnD(gameLogic_io_btnD),
    .io_songInput(gameLogic_io_songInput),
    .io_songStop(gameLogic_io_songStop),
    .io_spriteXPosition_0(gameLogic_io_spriteXPosition_0),
    .io_spriteYPosition_0(gameLogic_io_spriteYPosition_0),
    .io_spriteFlipHorizontal_0(gameLogic_io_spriteFlipHorizontal_0),
    .io_newFrame(gameLogic_io_newFrame),
    .io_frameUpdateDone(gameLogic_io_frameUpdateDone)
  );
  assign io_vgaRed = graphicEngineVGA_io_vgaRed; // @[GameTop.scala 104:13]
  assign io_vgaBlue = graphicEngineVGA_io_vgaBlue; // @[GameTop.scala 106:14]
  assign io_vgaGreen = graphicEngineVGA_io_vgaGreen; // @[GameTop.scala 105:15]
  assign io_Hsync = graphicEngineVGA_io_Hsync; // @[GameTop.scala 107:12]
  assign io_Vsync = graphicEngineVGA_io_Vsync; // @[GameTop.scala 108:12]
  assign io_soundOutput_0 = soundEngine_io_output_0; // @[GameTop.scala 122:18]
  assign io_missingFrameError = graphicEngineVGA_io_missingFrameError; // @[GameTop.scala 125:24]
  assign graphicEngineVGA_clock = clock;
  assign graphicEngineVGA_reset = _T_3 ? 1'h0 : 1'h1; // @[GameTop.scala 88:26]
  assign graphicEngineVGA_io_spriteXPosition_0 = gameLogic_io_spriteXPosition_0; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_0 = gameLogic_io_spriteYPosition_0; // @[GameTop.scala 131:39]
  assign graphicEngineVGA_io_spriteFlipHorizontal_0 = gameLogic_io_spriteFlipHorizontal_0; // @[GameTop.scala 133:44]
  assign graphicEngineVGA_io_frameUpdateDone = gameLogic_io_frameUpdateDone; // @[GameTop.scala 154:39]
  assign soundEngine_clock = clock;
  assign soundEngine_reset = reset;
  assign soundEngine_io_input = gameLogic_io_songInput; // @[GameTop.scala 119:24]
  assign soundEngine_io_stop = gameLogic_io_songStop; // @[GameTop.scala 120:23]
  assign gameLogic_clock = clock;
  assign gameLogic_reset = _T_3 ? 1'h0 : 1'h1; // @[GameTop.scala 89:19]
  assign gameLogic_io_btnC = btnCState; // @[GameTop.scala 97:21]
  assign gameLogic_io_btnU = btnUState; // @[GameTop.scala 98:21]
  assign gameLogic_io_btnL = btnLState; // @[GameTop.scala 99:21]
  assign gameLogic_io_btnR = btnRState; // @[GameTop.scala 100:21]
  assign gameLogic_io_btnD = btnDState; // @[GameTop.scala 101:21]
  assign gameLogic_io_newFrame = graphicEngineVGA_io_newFrame; // @[GameTop.scala 153:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounceCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  resetReleaseCounter = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  _T_7_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_7_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_7_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btnCState = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_9_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_9_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_9_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btnUState = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_11_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_11_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_11_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btnLState = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_13_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_13_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_13_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btnRState = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_15_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_15_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_15_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  btnDState = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      debounceCounter <= 21'h0;
    end else if (debounceSampleEn) begin
      debounceCounter <= 21'h0;
    end else begin
      debounceCounter <= _T_2;
    end
    if (reset) begin
      resetReleaseCounter <= 22'h0;
    end else if (!(_T_3)) begin
      resetReleaseCounter <= _T_5;
    end
    if (reset) begin
      _T_7_0 <= 1'h0;
    end else begin
      _T_7_0 <= _T_7_1;
    end
    if (reset) begin
      _T_7_1 <= 1'h0;
    end else begin
      _T_7_1 <= _T_7_2;
    end
    if (reset) begin
      _T_7_2 <= 1'h0;
    end else begin
      _T_7_2 <= io_btnC;
    end
    if (reset) begin
      btnCState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnCState <= _T_7_0;
    end
    if (reset) begin
      _T_9_0 <= 1'h0;
    end else begin
      _T_9_0 <= _T_9_1;
    end
    if (reset) begin
      _T_9_1 <= 1'h0;
    end else begin
      _T_9_1 <= _T_9_2;
    end
    if (reset) begin
      _T_9_2 <= 1'h0;
    end else begin
      _T_9_2 <= io_btnU;
    end
    if (reset) begin
      btnUState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnUState <= _T_9_0;
    end
    if (reset) begin
      _T_11_0 <= 1'h0;
    end else begin
      _T_11_0 <= _T_11_1;
    end
    if (reset) begin
      _T_11_1 <= 1'h0;
    end else begin
      _T_11_1 <= _T_11_2;
    end
    if (reset) begin
      _T_11_2 <= 1'h0;
    end else begin
      _T_11_2 <= io_btnL;
    end
    if (reset) begin
      btnLState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnLState <= _T_11_0;
    end
    if (reset) begin
      _T_13_0 <= 1'h0;
    end else begin
      _T_13_0 <= _T_13_1;
    end
    if (reset) begin
      _T_13_1 <= 1'h0;
    end else begin
      _T_13_1 <= _T_13_2;
    end
    if (reset) begin
      _T_13_2 <= 1'h0;
    end else begin
      _T_13_2 <= io_btnR;
    end
    if (reset) begin
      btnRState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnRState <= _T_13_0;
    end
    if (reset) begin
      _T_15_0 <= 1'h0;
    end else begin
      _T_15_0 <= _T_15_1;
    end
    if (reset) begin
      _T_15_1 <= 1'h0;
    end else begin
      _T_15_1 <= _T_15_2;
    end
    if (reset) begin
      _T_15_2 <= 1'h0;
    end else begin
      _T_15_2 <= io_btnD;
    end
    if (reset) begin
      btnDState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnDState <= _T_15_0;
    end
  end
endmodule
module Top(
  input        clock,
  input        reset,
  input        io_btnC,
  input        io_btnU,
  input        io_btnL,
  input        io_btnR,
  input        io_btnD,
  output [3:0] io_vgaRed,
  output [3:0] io_vgaGreen,
  output [3:0] io_vgaBlue,
  output       io_Hsync,
  output       io_Vsync,
  input        io_sw_0,
  input        io_sw_1,
  input        io_sw_2,
  input        io_sw_3,
  input        io_sw_4,
  input        io_sw_5,
  input        io_sw_6,
  input        io_sw_7,
  output       io_led_0,
  output       io_led_1,
  output       io_led_2,
  output       io_led_3,
  output       io_led_4,
  output       io_led_5,
  output       io_led_6,
  output       io_led_7,
  output       io_soundOutput_0,
  output       io_missingFrameError,
  output       io_backBufferWriteError,
  output       io_viewBoxOutOfRangeError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  gameTop_clock; // @[Top.scala 44:23]
  wire  gameTop_reset; // @[Top.scala 44:23]
  wire  gameTop_io_btnC; // @[Top.scala 44:23]
  wire  gameTop_io_btnU; // @[Top.scala 44:23]
  wire  gameTop_io_btnL; // @[Top.scala 44:23]
  wire  gameTop_io_btnR; // @[Top.scala 44:23]
  wire  gameTop_io_btnD; // @[Top.scala 44:23]
  wire [3:0] gameTop_io_vgaRed; // @[Top.scala 44:23]
  wire [3:0] gameTop_io_vgaBlue; // @[Top.scala 44:23]
  wire [3:0] gameTop_io_vgaGreen; // @[Top.scala 44:23]
  wire  gameTop_io_Hsync; // @[Top.scala 44:23]
  wire  gameTop_io_Vsync; // @[Top.scala 44:23]
  wire  gameTop_io_soundOutput_0; // @[Top.scala 44:23]
  wire  gameTop_io_missingFrameError; // @[Top.scala 44:23]
  reg  _T_1; // @[Top.scala 49:48]
  reg  _T_2; // @[Top.scala 49:40]
  reg  _T_3; // @[Top.scala 49:32]
  reg  pipeResetReg_0; // @[Top.scala 54:25]
  reg  pipeResetReg_1; // @[Top.scala 54:25]
  reg  pipeResetReg_2; // @[Top.scala 54:25]
  reg  pipeResetReg_3; // @[Top.scala 54:25]
  reg  pipeResetReg_4; // @[Top.scala 54:25]
  wire [4:0] _T_7 = {pipeResetReg_4,pipeResetReg_3,pipeResetReg_2,pipeResetReg_1,pipeResetReg_0}; // @[Top.scala 59:33]
  GameTop gameTop ( // @[Top.scala 44:23]
    .clock(gameTop_clock),
    .reset(gameTop_reset),
    .io_btnC(gameTop_io_btnC),
    .io_btnU(gameTop_io_btnU),
    .io_btnL(gameTop_io_btnL),
    .io_btnR(gameTop_io_btnR),
    .io_btnD(gameTop_io_btnD),
    .io_vgaRed(gameTop_io_vgaRed),
    .io_vgaBlue(gameTop_io_vgaBlue),
    .io_vgaGreen(gameTop_io_vgaGreen),
    .io_Hsync(gameTop_io_Hsync),
    .io_Vsync(gameTop_io_Vsync),
    .io_soundOutput_0(gameTop_io_soundOutput_0),
    .io_missingFrameError(gameTop_io_missingFrameError)
  );
  assign io_vgaRed = gameTop_io_vgaRed; // @[Top.scala 62:14]
  assign io_vgaGreen = gameTop_io_vgaGreen; // @[Top.scala 62:14]
  assign io_vgaBlue = gameTop_io_vgaBlue; // @[Top.scala 62:14]
  assign io_Hsync = gameTop_io_Hsync; // @[Top.scala 62:14]
  assign io_Vsync = gameTop_io_Vsync; // @[Top.scala 62:14]
  assign io_led_0 = 1'h0; // @[Top.scala 62:14]
  assign io_led_1 = 1'h0; // @[Top.scala 62:14]
  assign io_led_2 = 1'h0; // @[Top.scala 62:14]
  assign io_led_3 = 1'h0; // @[Top.scala 62:14]
  assign io_led_4 = 1'h0; // @[Top.scala 62:14]
  assign io_led_5 = 1'h0; // @[Top.scala 62:14]
  assign io_led_6 = 1'h0; // @[Top.scala 62:14]
  assign io_led_7 = 1'h0; // @[Top.scala 62:14]
  assign io_soundOutput_0 = gameTop_io_soundOutput_0; // @[Top.scala 62:14]
  assign io_missingFrameError = gameTop_io_missingFrameError; // @[Top.scala 62:14]
  assign io_backBufferWriteError = 1'h0; // @[Top.scala 62:14]
  assign io_viewBoxOutOfRangeError = 1'h0; // @[Top.scala 62:14]
  assign gameTop_clock = clock;
  assign gameTop_reset = |_T_7; // @[Top.scala 59:17]
  assign gameTop_io_btnC = io_btnC; // @[Top.scala 62:14]
  assign gameTop_io_btnU = io_btnU; // @[Top.scala 62:14]
  assign gameTop_io_btnL = io_btnL; // @[Top.scala 62:14]
  assign gameTop_io_btnR = io_btnR; // @[Top.scala 62:14]
  assign gameTop_io_btnD = io_btnD; // @[Top.scala 62:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_2 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipeResetReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipeResetReg_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pipeResetReg_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipeResetReg_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pipeResetReg_4 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= reset;
    _T_2 <= _T_1;
    _T_3 <= _T_2;
    pipeResetReg_0 <= pipeResetReg_1;
    pipeResetReg_1 <= pipeResetReg_2;
    pipeResetReg_2 <= pipeResetReg_3;
    pipeResetReg_3 <= pipeResetReg_4;
    pipeResetReg_4 <= ~_T_3;
  end
endmodule
