module Memory(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_1(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_2(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_3(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_4(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_5(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_6(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_7(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_8(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_8.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_9(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_9.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_10(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_10.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_11(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_11.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_12(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_12.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_13(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_13.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_14(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_14.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_15(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_15.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_16(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_16.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_17(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_17.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_18(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_18.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_19(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_19.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_20(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_20.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_21(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_21.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_22(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_22.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_23(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_23.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_24(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_24.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_25(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_25.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_26(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_26.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_27(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_27.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_28(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_28.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_29(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_29.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_30(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_30.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_31(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/backtile_init_31.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_64(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead,
  input         io_writeEnable,
  input  [4:0]  io_dataWrite
);
  wire  RamSpWf_clk; // @[Memory.scala 57:26]
  wire  RamSpWf_we; // @[Memory.scala 57:26]
  wire  RamSpWf_en; // @[Memory.scala 57:26]
  wire [10:0] RamSpWf_addr; // @[Memory.scala 57:26]
  wire [4:0] RamSpWf_di; // @[Memory.scala 57:26]
  wire [4:0] RamSpWf_dout; // @[Memory.scala 57:26]
  RamSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5)) RamSpWf ( // @[Memory.scala 57:26]
    .clk(RamSpWf_clk),
    .we(RamSpWf_we),
    .en(RamSpWf_en),
    .addr(RamSpWf_addr),
    .di(RamSpWf_di),
    .dout(RamSpWf_dout)
  );
  assign io_dataRead = RamSpWf_dout; // @[Memory.scala 63:17]
  assign RamSpWf_clk = clock; // @[Memory.scala 58:21]
  assign RamSpWf_we = io_writeEnable; // @[Memory.scala 59:20]
  assign RamSpWf_en = 1'h1; // @[Memory.scala 60:20]
  assign RamSpWf_addr = io_address; // @[Memory.scala 61:22]
  assign RamSpWf_di = io_dataWrite; // @[Memory.scala 62:20]
endmodule
module Memory_68(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [10:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5), .LOAD_FILE("memory_init/backbuffer_init0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 5'h0; // @[Memory.scala 70:20]
endmodule
module Memory_69(
  input         clock,
  input  [10:0] io_address,
  output [4:0]  io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [10:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [4:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(11), .DATA_WIDTH(5), .LOAD_FILE("memory_init/backbuffer_init1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 5'h0; // @[Memory.scala 70:20]
endmodule
module Memory_70(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_71(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_72(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_73(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_74(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_75(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_76(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_77(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_78(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_8.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_79(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_9.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_80(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_10.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_81(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_11.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_82(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_12.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_83(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_13.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_84(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_14.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_85(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_15.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_86(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_16.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_87(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_17.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_88(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_18.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_89(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_19.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_90(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_20.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_91(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_21.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_92(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_22.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_93(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_23.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_94(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_24.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_95(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_25.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_96(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_26.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_97(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_27.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_98(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_28.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_99(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_29.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_100(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_30.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_101(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_31.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_102(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_32.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_103(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_33.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_104(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_34.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_105(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_35.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_106(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_36.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_107(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_37.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_108(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_38.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_109(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_39.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_110(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_40.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_111(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_41.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_112(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_42.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_113(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_43.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_114(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_44.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_115(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_45.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_116(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_46.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_117(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_47.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_118(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_48.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_119(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_49.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_120(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_50.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_121(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_51.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_122(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_52.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_123(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_53.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_124(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_54.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_125(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_55.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_126(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_56.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_127(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_57.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_128(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_58.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_129(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_59.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_130(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_60.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_131(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_61.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_132(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_62.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_133(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_63.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_134(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_64.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_135(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_65.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_136(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_66.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_137(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_67.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_138(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_68.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_139(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_69.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_140(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_70.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_141(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_71.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_142(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_72.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_143(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_73.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_144(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_74.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_145(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_75.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_146(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_76.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_147(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_77.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_148(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_78.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_149(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_79.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_150(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_80.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_151(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_81.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_152(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_82.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_153(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_83.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_154(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_84.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_155(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_85.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_156(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_86.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_157(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_87.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_158(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_88.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_159(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_89.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_160(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_90.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_161(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_91.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_162(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_92.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_163(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_93.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_164(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_94.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_165(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_95.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_166(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_96.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_167(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_97.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_168(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_98.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_169(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_99.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_170(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_100.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_171(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_101.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_172(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_102.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_173(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_103.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_174(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_104.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_175(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_105.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_176(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_106.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_177(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_107.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_178(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_108.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_179(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_109.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_180(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_110.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_181(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_111.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_182(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_112.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_183(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_113.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_184(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_114.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_185(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_115.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_186(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_116.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_187(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_117.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_188(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_118.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_189(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_119.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_190(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_120.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_191(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_121.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_192(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_122.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_193(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_123.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_194(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_124.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_195(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_125.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_196(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_126.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module Memory_197(
  input        clock,
  input  [9:0] io_address,
  output [6:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [9:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [6:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(10), .DATA_WIDTH(7), .LOAD_FILE("memory_init/sprite_init_127.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 7'h0; // @[Memory.scala 70:20]
endmodule
module MultiHotPriortyReductionTree(
  input  [5:0] io_dataInput_0,
  input  [5:0] io_dataInput_1,
  input  [5:0] io_dataInput_2,
  input  [5:0] io_dataInput_3,
  input  [5:0] io_dataInput_4,
  input  [5:0] io_dataInput_5,
  input  [5:0] io_dataInput_6,
  input  [5:0] io_dataInput_7,
  input  [5:0] io_dataInput_8,
  input  [5:0] io_dataInput_9,
  input  [5:0] io_dataInput_10,
  input  [5:0] io_dataInput_11,
  input  [5:0] io_dataInput_12,
  input  [5:0] io_dataInput_13,
  input  [5:0] io_dataInput_14,
  input  [5:0] io_dataInput_15,
  input  [5:0] io_dataInput_16,
  input  [5:0] io_dataInput_17,
  input  [5:0] io_dataInput_18,
  input  [5:0] io_dataInput_19,
  input  [5:0] io_dataInput_20,
  input  [5:0] io_dataInput_21,
  input  [5:0] io_dataInput_22,
  input  [5:0] io_dataInput_23,
  input  [5:0] io_dataInput_24,
  input  [5:0] io_dataInput_25,
  input  [5:0] io_dataInput_26,
  input  [5:0] io_dataInput_27,
  input  [5:0] io_dataInput_28,
  input  [5:0] io_dataInput_29,
  input  [5:0] io_dataInput_30,
  input  [5:0] io_dataInput_31,
  input  [5:0] io_dataInput_32,
  input  [5:0] io_dataInput_33,
  input  [5:0] io_dataInput_34,
  input  [5:0] io_dataInput_35,
  input  [5:0] io_dataInput_36,
  input  [5:0] io_dataInput_37,
  input  [5:0] io_dataInput_38,
  input  [5:0] io_dataInput_39,
  input  [5:0] io_dataInput_40,
  input  [5:0] io_dataInput_41,
  input  [5:0] io_dataInput_42,
  input  [5:0] io_dataInput_43,
  input  [5:0] io_dataInput_44,
  input  [5:0] io_dataInput_45,
  input  [5:0] io_dataInput_46,
  input  [5:0] io_dataInput_47,
  input  [5:0] io_dataInput_48,
  input  [5:0] io_dataInput_49,
  input  [5:0] io_dataInput_50,
  input  [5:0] io_dataInput_51,
  input  [5:0] io_dataInput_52,
  input  [5:0] io_dataInput_53,
  input  [5:0] io_dataInput_54,
  input  [5:0] io_dataInput_55,
  input  [5:0] io_dataInput_56,
  input  [5:0] io_dataInput_57,
  input  [5:0] io_dataInput_58,
  input  [5:0] io_dataInput_59,
  input  [5:0] io_dataInput_60,
  input  [5:0] io_dataInput_61,
  input  [5:0] io_dataInput_62,
  input  [5:0] io_dataInput_63,
  input  [5:0] io_dataInput_64,
  input  [5:0] io_dataInput_65,
  input  [5:0] io_dataInput_66,
  input  [5:0] io_dataInput_67,
  input  [5:0] io_dataInput_68,
  input  [5:0] io_dataInput_69,
  input  [5:0] io_dataInput_70,
  input  [5:0] io_dataInput_71,
  input  [5:0] io_dataInput_72,
  input  [5:0] io_dataInput_73,
  input  [5:0] io_dataInput_74,
  input  [5:0] io_dataInput_75,
  input  [5:0] io_dataInput_76,
  input  [5:0] io_dataInput_77,
  input  [5:0] io_dataInput_78,
  input  [5:0] io_dataInput_79,
  input  [5:0] io_dataInput_80,
  input  [5:0] io_dataInput_81,
  input  [5:0] io_dataInput_82,
  input  [5:0] io_dataInput_83,
  input  [5:0] io_dataInput_84,
  input  [5:0] io_dataInput_85,
  input  [5:0] io_dataInput_86,
  input  [5:0] io_dataInput_87,
  input  [5:0] io_dataInput_88,
  input  [5:0] io_dataInput_89,
  input  [5:0] io_dataInput_90,
  input  [5:0] io_dataInput_91,
  input  [5:0] io_dataInput_92,
  input  [5:0] io_dataInput_93,
  input  [5:0] io_dataInput_94,
  input  [5:0] io_dataInput_95,
  input  [5:0] io_dataInput_96,
  input  [5:0] io_dataInput_97,
  input  [5:0] io_dataInput_98,
  input  [5:0] io_dataInput_99,
  input  [5:0] io_dataInput_100,
  input  [5:0] io_dataInput_101,
  input  [5:0] io_dataInput_102,
  input  [5:0] io_dataInput_103,
  input  [5:0] io_dataInput_104,
  input  [5:0] io_dataInput_105,
  input  [5:0] io_dataInput_106,
  input  [5:0] io_dataInput_107,
  input  [5:0] io_dataInput_108,
  input  [5:0] io_dataInput_109,
  input  [5:0] io_dataInput_110,
  input  [5:0] io_dataInput_111,
  input  [5:0] io_dataInput_112,
  input  [5:0] io_dataInput_113,
  input  [5:0] io_dataInput_114,
  input  [5:0] io_dataInput_115,
  input  [5:0] io_dataInput_116,
  input  [5:0] io_dataInput_117,
  input  [5:0] io_dataInput_118,
  input  [5:0] io_dataInput_119,
  input  [5:0] io_dataInput_120,
  input  [5:0] io_dataInput_121,
  input  [5:0] io_dataInput_122,
  input  [5:0] io_dataInput_123,
  input  [5:0] io_dataInput_124,
  input  [5:0] io_dataInput_125,
  input  [5:0] io_dataInput_126,
  input  [5:0] io_dataInput_127,
  input        io_selectInput_0,
  input        io_selectInput_1,
  input        io_selectInput_2,
  input        io_selectInput_3,
  input        io_selectInput_4,
  input        io_selectInput_5,
  input        io_selectInput_6,
  input        io_selectInput_7,
  input        io_selectInput_8,
  input        io_selectInput_9,
  input        io_selectInput_10,
  input        io_selectInput_11,
  input        io_selectInput_12,
  input        io_selectInput_13,
  input        io_selectInput_14,
  input        io_selectInput_15,
  input        io_selectInput_16,
  input        io_selectInput_17,
  input        io_selectInput_18,
  input        io_selectInput_19,
  input        io_selectInput_20,
  input        io_selectInput_21,
  input        io_selectInput_22,
  input        io_selectInput_23,
  input        io_selectInput_24,
  input        io_selectInput_25,
  input        io_selectInput_26,
  input        io_selectInput_27,
  input        io_selectInput_28,
  input        io_selectInput_29,
  input        io_selectInput_30,
  input        io_selectInput_31,
  input        io_selectInput_32,
  input        io_selectInput_33,
  input        io_selectInput_34,
  input        io_selectInput_35,
  input        io_selectInput_36,
  input        io_selectInput_37,
  input        io_selectInput_38,
  input        io_selectInput_39,
  input        io_selectInput_40,
  input        io_selectInput_41,
  input        io_selectInput_42,
  input        io_selectInput_43,
  input        io_selectInput_44,
  input        io_selectInput_45,
  input        io_selectInput_46,
  input        io_selectInput_47,
  input        io_selectInput_48,
  input        io_selectInput_49,
  input        io_selectInput_50,
  input        io_selectInput_51,
  input        io_selectInput_52,
  input        io_selectInput_53,
  input        io_selectInput_54,
  input        io_selectInput_55,
  input        io_selectInput_56,
  input        io_selectInput_57,
  input        io_selectInput_58,
  input        io_selectInput_59,
  input        io_selectInput_60,
  input        io_selectInput_61,
  input        io_selectInput_62,
  input        io_selectInput_63,
  input        io_selectInput_64,
  input        io_selectInput_65,
  input        io_selectInput_66,
  input        io_selectInput_67,
  input        io_selectInput_68,
  input        io_selectInput_69,
  input        io_selectInput_70,
  input        io_selectInput_71,
  input        io_selectInput_72,
  input        io_selectInput_73,
  input        io_selectInput_74,
  input        io_selectInput_75,
  input        io_selectInput_76,
  input        io_selectInput_77,
  input        io_selectInput_78,
  input        io_selectInput_79,
  input        io_selectInput_80,
  input        io_selectInput_81,
  input        io_selectInput_82,
  input        io_selectInput_83,
  input        io_selectInput_84,
  input        io_selectInput_85,
  input        io_selectInput_86,
  input        io_selectInput_87,
  input        io_selectInput_88,
  input        io_selectInput_89,
  input        io_selectInput_90,
  input        io_selectInput_91,
  input        io_selectInput_92,
  input        io_selectInput_93,
  input        io_selectInput_94,
  input        io_selectInput_95,
  input        io_selectInput_96,
  input        io_selectInput_97,
  input        io_selectInput_98,
  input        io_selectInput_99,
  input        io_selectInput_100,
  input        io_selectInput_101,
  input        io_selectInput_102,
  input        io_selectInput_103,
  input        io_selectInput_104,
  input        io_selectInput_105,
  input        io_selectInput_106,
  input        io_selectInput_107,
  input        io_selectInput_108,
  input        io_selectInput_109,
  input        io_selectInput_110,
  input        io_selectInput_111,
  input        io_selectInput_112,
  input        io_selectInput_113,
  input        io_selectInput_114,
  input        io_selectInput_115,
  input        io_selectInput_116,
  input        io_selectInput_117,
  input        io_selectInput_118,
  input        io_selectInput_119,
  input        io_selectInput_120,
  input        io_selectInput_121,
  input        io_selectInput_122,
  input        io_selectInput_123,
  input        io_selectInput_124,
  input        io_selectInput_125,
  input        io_selectInput_126,
  input        io_selectInput_127,
  output [5:0] io_dataOutput,
  output       io_selectOutput
);
  wire  selectNodeOutputs_63 = io_selectInput_0 | io_selectInput_1; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_64 = io_selectInput_2 | io_selectInput_3; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_31 = selectNodeOutputs_63 | selectNodeOutputs_64; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_65 = io_selectInput_4 | io_selectInput_5; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_66 = io_selectInput_6 | io_selectInput_7; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_32 = selectNodeOutputs_65 | selectNodeOutputs_66; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_15 = selectNodeOutputs_31 | selectNodeOutputs_32; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_67 = io_selectInput_8 | io_selectInput_9; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_68 = io_selectInput_10 | io_selectInput_11; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_33 = selectNodeOutputs_67 | selectNodeOutputs_68; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_69 = io_selectInput_12 | io_selectInput_13; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_70 = io_selectInput_14 | io_selectInput_15; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_34 = selectNodeOutputs_69 | selectNodeOutputs_70; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_16 = selectNodeOutputs_33 | selectNodeOutputs_34; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_7 = selectNodeOutputs_15 | selectNodeOutputs_16; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_71 = io_selectInput_16 | io_selectInput_17; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_72 = io_selectInput_18 | io_selectInput_19; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_35 = selectNodeOutputs_71 | selectNodeOutputs_72; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_73 = io_selectInput_20 | io_selectInput_21; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_74 = io_selectInput_22 | io_selectInput_23; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_36 = selectNodeOutputs_73 | selectNodeOutputs_74; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_17 = selectNodeOutputs_35 | selectNodeOutputs_36; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_75 = io_selectInput_24 | io_selectInput_25; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_76 = io_selectInput_26 | io_selectInput_27; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_37 = selectNodeOutputs_75 | selectNodeOutputs_76; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_77 = io_selectInput_28 | io_selectInput_29; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_78 = io_selectInput_30 | io_selectInput_31; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_38 = selectNodeOutputs_77 | selectNodeOutputs_78; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_18 = selectNodeOutputs_37 | selectNodeOutputs_38; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_8 = selectNodeOutputs_17 | selectNodeOutputs_18; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_3 = selectNodeOutputs_7 | selectNodeOutputs_8; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_79 = io_selectInput_32 | io_selectInput_33; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_80 = io_selectInput_34 | io_selectInput_35; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_39 = selectNodeOutputs_79 | selectNodeOutputs_80; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_81 = io_selectInput_36 | io_selectInput_37; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_82 = io_selectInput_38 | io_selectInput_39; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_40 = selectNodeOutputs_81 | selectNodeOutputs_82; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_19 = selectNodeOutputs_39 | selectNodeOutputs_40; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_83 = io_selectInput_40 | io_selectInput_41; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_84 = io_selectInput_42 | io_selectInput_43; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_41 = selectNodeOutputs_83 | selectNodeOutputs_84; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_85 = io_selectInput_44 | io_selectInput_45; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_86 = io_selectInput_46 | io_selectInput_47; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_42 = selectNodeOutputs_85 | selectNodeOutputs_86; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_20 = selectNodeOutputs_41 | selectNodeOutputs_42; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_9 = selectNodeOutputs_19 | selectNodeOutputs_20; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_87 = io_selectInput_48 | io_selectInput_49; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_88 = io_selectInput_50 | io_selectInput_51; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_43 = selectNodeOutputs_87 | selectNodeOutputs_88; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_89 = io_selectInput_52 | io_selectInput_53; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_90 = io_selectInput_54 | io_selectInput_55; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_44 = selectNodeOutputs_89 | selectNodeOutputs_90; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_21 = selectNodeOutputs_43 | selectNodeOutputs_44; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_91 = io_selectInput_56 | io_selectInput_57; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_92 = io_selectInput_58 | io_selectInput_59; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_45 = selectNodeOutputs_91 | selectNodeOutputs_92; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_93 = io_selectInput_60 | io_selectInput_61; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_94 = io_selectInput_62 | io_selectInput_63; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_46 = selectNodeOutputs_93 | selectNodeOutputs_94; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_22 = selectNodeOutputs_45 | selectNodeOutputs_46; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_10 = selectNodeOutputs_21 | selectNodeOutputs_22; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_4 = selectNodeOutputs_9 | selectNodeOutputs_10; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_1 = selectNodeOutputs_3 | selectNodeOutputs_4; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_63 = io_selectInput_0 ? io_dataInput_0 : io_dataInput_1; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_64 = io_selectInput_2 ? io_dataInput_2 : io_dataInput_3; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_31 = selectNodeOutputs_63 ? dataNodeOutputs_63 : dataNodeOutputs_64; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_65 = io_selectInput_4 ? io_dataInput_4 : io_dataInput_5; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_66 = io_selectInput_6 ? io_dataInput_6 : io_dataInput_7; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_32 = selectNodeOutputs_65 ? dataNodeOutputs_65 : dataNodeOutputs_66; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_15 = selectNodeOutputs_31 ? dataNodeOutputs_31 : dataNodeOutputs_32; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_67 = io_selectInput_8 ? io_dataInput_8 : io_dataInput_9; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_68 = io_selectInput_10 ? io_dataInput_10 : io_dataInput_11; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_33 = selectNodeOutputs_67 ? dataNodeOutputs_67 : dataNodeOutputs_68; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_69 = io_selectInput_12 ? io_dataInput_12 : io_dataInput_13; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_70 = io_selectInput_14 ? io_dataInput_14 : io_dataInput_15; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_34 = selectNodeOutputs_69 ? dataNodeOutputs_69 : dataNodeOutputs_70; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_16 = selectNodeOutputs_33 ? dataNodeOutputs_33 : dataNodeOutputs_34; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_7 = selectNodeOutputs_15 ? dataNodeOutputs_15 : dataNodeOutputs_16; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_71 = io_selectInput_16 ? io_dataInput_16 : io_dataInput_17; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_72 = io_selectInput_18 ? io_dataInput_18 : io_dataInput_19; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_35 = selectNodeOutputs_71 ? dataNodeOutputs_71 : dataNodeOutputs_72; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_73 = io_selectInput_20 ? io_dataInput_20 : io_dataInput_21; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_74 = io_selectInput_22 ? io_dataInput_22 : io_dataInput_23; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_36 = selectNodeOutputs_73 ? dataNodeOutputs_73 : dataNodeOutputs_74; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_17 = selectNodeOutputs_35 ? dataNodeOutputs_35 : dataNodeOutputs_36; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_75 = io_selectInput_24 ? io_dataInput_24 : io_dataInput_25; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_76 = io_selectInput_26 ? io_dataInput_26 : io_dataInput_27; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_37 = selectNodeOutputs_75 ? dataNodeOutputs_75 : dataNodeOutputs_76; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_77 = io_selectInput_28 ? io_dataInput_28 : io_dataInput_29; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_78 = io_selectInput_30 ? io_dataInput_30 : io_dataInput_31; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_38 = selectNodeOutputs_77 ? dataNodeOutputs_77 : dataNodeOutputs_78; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_18 = selectNodeOutputs_37 ? dataNodeOutputs_37 : dataNodeOutputs_38; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_8 = selectNodeOutputs_17 ? dataNodeOutputs_17 : dataNodeOutputs_18; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_3 = selectNodeOutputs_7 ? dataNodeOutputs_7 : dataNodeOutputs_8; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_79 = io_selectInput_32 ? io_dataInput_32 : io_dataInput_33; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_80 = io_selectInput_34 ? io_dataInput_34 : io_dataInput_35; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_39 = selectNodeOutputs_79 ? dataNodeOutputs_79 : dataNodeOutputs_80; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_81 = io_selectInput_36 ? io_dataInput_36 : io_dataInput_37; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_82 = io_selectInput_38 ? io_dataInput_38 : io_dataInput_39; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_40 = selectNodeOutputs_81 ? dataNodeOutputs_81 : dataNodeOutputs_82; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_19 = selectNodeOutputs_39 ? dataNodeOutputs_39 : dataNodeOutputs_40; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_83 = io_selectInput_40 ? io_dataInput_40 : io_dataInput_41; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_84 = io_selectInput_42 ? io_dataInput_42 : io_dataInput_43; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_41 = selectNodeOutputs_83 ? dataNodeOutputs_83 : dataNodeOutputs_84; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_85 = io_selectInput_44 ? io_dataInput_44 : io_dataInput_45; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_86 = io_selectInput_46 ? io_dataInput_46 : io_dataInput_47; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_42 = selectNodeOutputs_85 ? dataNodeOutputs_85 : dataNodeOutputs_86; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_20 = selectNodeOutputs_41 ? dataNodeOutputs_41 : dataNodeOutputs_42; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_9 = selectNodeOutputs_19 ? dataNodeOutputs_19 : dataNodeOutputs_20; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_87 = io_selectInput_48 ? io_dataInput_48 : io_dataInput_49; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_88 = io_selectInput_50 ? io_dataInput_50 : io_dataInput_51; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_43 = selectNodeOutputs_87 ? dataNodeOutputs_87 : dataNodeOutputs_88; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_89 = io_selectInput_52 ? io_dataInput_52 : io_dataInput_53; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_90 = io_selectInput_54 ? io_dataInput_54 : io_dataInput_55; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_44 = selectNodeOutputs_89 ? dataNodeOutputs_89 : dataNodeOutputs_90; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_21 = selectNodeOutputs_43 ? dataNodeOutputs_43 : dataNodeOutputs_44; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_91 = io_selectInput_56 ? io_dataInput_56 : io_dataInput_57; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_92 = io_selectInput_58 ? io_dataInput_58 : io_dataInput_59; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_45 = selectNodeOutputs_91 ? dataNodeOutputs_91 : dataNodeOutputs_92; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_93 = io_selectInput_60 ? io_dataInput_60 : io_dataInput_61; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_94 = io_selectInput_62 ? io_dataInput_62 : io_dataInput_63; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_46 = selectNodeOutputs_93 ? dataNodeOutputs_93 : dataNodeOutputs_94; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_22 = selectNodeOutputs_45 ? dataNodeOutputs_45 : dataNodeOutputs_46; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_10 = selectNodeOutputs_21 ? dataNodeOutputs_21 : dataNodeOutputs_22; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_4 = selectNodeOutputs_9 ? dataNodeOutputs_9 : dataNodeOutputs_10; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_1 = selectNodeOutputs_3 ? dataNodeOutputs_3 : dataNodeOutputs_4; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_95 = io_selectInput_64 | io_selectInput_65; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_96 = io_selectInput_66 | io_selectInput_67; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_47 = selectNodeOutputs_95 | selectNodeOutputs_96; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_97 = io_selectInput_68 | io_selectInput_69; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_98 = io_selectInput_70 | io_selectInput_71; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_48 = selectNodeOutputs_97 | selectNodeOutputs_98; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_23 = selectNodeOutputs_47 | selectNodeOutputs_48; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_99 = io_selectInput_72 | io_selectInput_73; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_100 = io_selectInput_74 | io_selectInput_75; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_49 = selectNodeOutputs_99 | selectNodeOutputs_100; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_101 = io_selectInput_76 | io_selectInput_77; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_102 = io_selectInput_78 | io_selectInput_79; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_50 = selectNodeOutputs_101 | selectNodeOutputs_102; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_24 = selectNodeOutputs_49 | selectNodeOutputs_50; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_11 = selectNodeOutputs_23 | selectNodeOutputs_24; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_103 = io_selectInput_80 | io_selectInput_81; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_104 = io_selectInput_82 | io_selectInput_83; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_51 = selectNodeOutputs_103 | selectNodeOutputs_104; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_105 = io_selectInput_84 | io_selectInput_85; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_106 = io_selectInput_86 | io_selectInput_87; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_52 = selectNodeOutputs_105 | selectNodeOutputs_106; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_25 = selectNodeOutputs_51 | selectNodeOutputs_52; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_107 = io_selectInput_88 | io_selectInput_89; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_108 = io_selectInput_90 | io_selectInput_91; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_53 = selectNodeOutputs_107 | selectNodeOutputs_108; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_109 = io_selectInput_92 | io_selectInput_93; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_110 = io_selectInput_94 | io_selectInput_95; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_54 = selectNodeOutputs_109 | selectNodeOutputs_110; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_26 = selectNodeOutputs_53 | selectNodeOutputs_54; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_12 = selectNodeOutputs_25 | selectNodeOutputs_26; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_5 = selectNodeOutputs_11 | selectNodeOutputs_12; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_95 = io_selectInput_64 ? io_dataInput_64 : io_dataInput_65; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_96 = io_selectInput_66 ? io_dataInput_66 : io_dataInput_67; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_47 = selectNodeOutputs_95 ? dataNodeOutputs_95 : dataNodeOutputs_96; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_97 = io_selectInput_68 ? io_dataInput_68 : io_dataInput_69; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_98 = io_selectInput_70 ? io_dataInput_70 : io_dataInput_71; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_48 = selectNodeOutputs_97 ? dataNodeOutputs_97 : dataNodeOutputs_98; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_23 = selectNodeOutputs_47 ? dataNodeOutputs_47 : dataNodeOutputs_48; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_99 = io_selectInput_72 ? io_dataInput_72 : io_dataInput_73; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_100 = io_selectInput_74 ? io_dataInput_74 : io_dataInput_75; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_49 = selectNodeOutputs_99 ? dataNodeOutputs_99 : dataNodeOutputs_100; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_101 = io_selectInput_76 ? io_dataInput_76 : io_dataInput_77; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_102 = io_selectInput_78 ? io_dataInput_78 : io_dataInput_79; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_50 = selectNodeOutputs_101 ? dataNodeOutputs_101 : dataNodeOutputs_102; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_24 = selectNodeOutputs_49 ? dataNodeOutputs_49 : dataNodeOutputs_50; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_11 = selectNodeOutputs_23 ? dataNodeOutputs_23 : dataNodeOutputs_24; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_103 = io_selectInput_80 ? io_dataInput_80 : io_dataInput_81; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_104 = io_selectInput_82 ? io_dataInput_82 : io_dataInput_83; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_51 = selectNodeOutputs_103 ? dataNodeOutputs_103 : dataNodeOutputs_104; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_105 = io_selectInput_84 ? io_dataInput_84 : io_dataInput_85; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_106 = io_selectInput_86 ? io_dataInput_86 : io_dataInput_87; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_52 = selectNodeOutputs_105 ? dataNodeOutputs_105 : dataNodeOutputs_106; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_25 = selectNodeOutputs_51 ? dataNodeOutputs_51 : dataNodeOutputs_52; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_107 = io_selectInput_88 ? io_dataInput_88 : io_dataInput_89; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_108 = io_selectInput_90 ? io_dataInput_90 : io_dataInput_91; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_53 = selectNodeOutputs_107 ? dataNodeOutputs_107 : dataNodeOutputs_108; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_109 = io_selectInput_92 ? io_dataInput_92 : io_dataInput_93; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_110 = io_selectInput_94 ? io_dataInput_94 : io_dataInput_95; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_54 = selectNodeOutputs_109 ? dataNodeOutputs_109 : dataNodeOutputs_110; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_26 = selectNodeOutputs_53 ? dataNodeOutputs_53 : dataNodeOutputs_54; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_12 = selectNodeOutputs_25 ? dataNodeOutputs_25 : dataNodeOutputs_26; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_5 = selectNodeOutputs_11 ? dataNodeOutputs_11 : dataNodeOutputs_12; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_111 = io_selectInput_96 | io_selectInput_97; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_112 = io_selectInput_98 | io_selectInput_99; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_55 = selectNodeOutputs_111 | selectNodeOutputs_112; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_113 = io_selectInput_100 | io_selectInput_101; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_114 = io_selectInput_102 | io_selectInput_103; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_56 = selectNodeOutputs_113 | selectNodeOutputs_114; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_27 = selectNodeOutputs_55 | selectNodeOutputs_56; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_115 = io_selectInput_104 | io_selectInput_105; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_116 = io_selectInput_106 | io_selectInput_107; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_57 = selectNodeOutputs_115 | selectNodeOutputs_116; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_117 = io_selectInput_108 | io_selectInput_109; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_118 = io_selectInput_110 | io_selectInput_111; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_58 = selectNodeOutputs_117 | selectNodeOutputs_118; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_28 = selectNodeOutputs_57 | selectNodeOutputs_58; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_13 = selectNodeOutputs_27 | selectNodeOutputs_28; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_111 = io_selectInput_96 ? io_dataInput_96 : io_dataInput_97; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_112 = io_selectInput_98 ? io_dataInput_98 : io_dataInput_99; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_55 = selectNodeOutputs_111 ? dataNodeOutputs_111 : dataNodeOutputs_112; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_113 = io_selectInput_100 ? io_dataInput_100 : io_dataInput_101; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_114 = io_selectInput_102 ? io_dataInput_102 : io_dataInput_103; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_56 = selectNodeOutputs_113 ? dataNodeOutputs_113 : dataNodeOutputs_114; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_27 = selectNodeOutputs_55 ? dataNodeOutputs_55 : dataNodeOutputs_56; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_115 = io_selectInput_104 ? io_dataInput_104 : io_dataInput_105; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_116 = io_selectInput_106 ? io_dataInput_106 : io_dataInput_107; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_57 = selectNodeOutputs_115 ? dataNodeOutputs_115 : dataNodeOutputs_116; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_117 = io_selectInput_108 ? io_dataInput_108 : io_dataInput_109; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_118 = io_selectInput_110 ? io_dataInput_110 : io_dataInput_111; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_58 = selectNodeOutputs_117 ? dataNodeOutputs_117 : dataNodeOutputs_118; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_28 = selectNodeOutputs_57 ? dataNodeOutputs_57 : dataNodeOutputs_58; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_13 = selectNodeOutputs_27 ? dataNodeOutputs_27 : dataNodeOutputs_28; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_119 = io_selectInput_112 | io_selectInput_113; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_120 = io_selectInput_114 | io_selectInput_115; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_59 = selectNodeOutputs_119 | selectNodeOutputs_120; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_121 = io_selectInput_116 | io_selectInput_117; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_122 = io_selectInput_118 | io_selectInput_119; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_60 = selectNodeOutputs_121 | selectNodeOutputs_122; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_29 = selectNodeOutputs_59 | selectNodeOutputs_60; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_119 = io_selectInput_112 ? io_dataInput_112 : io_dataInput_113; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_120 = io_selectInput_114 ? io_dataInput_114 : io_dataInput_115; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_59 = selectNodeOutputs_119 ? dataNodeOutputs_119 : dataNodeOutputs_120; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_121 = io_selectInput_116 ? io_dataInput_116 : io_dataInput_117; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_122 = io_selectInput_118 ? io_dataInput_118 : io_dataInput_119; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_60 = selectNodeOutputs_121 ? dataNodeOutputs_121 : dataNodeOutputs_122; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_29 = selectNodeOutputs_59 ? dataNodeOutputs_59 : dataNodeOutputs_60; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_123 = io_selectInput_120 | io_selectInput_121; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_124 = io_selectInput_122 | io_selectInput_123; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_61 = selectNodeOutputs_123 | selectNodeOutputs_124; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_123 = io_selectInput_120 ? io_dataInput_120 : io_dataInput_121; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_124 = io_selectInput_122 ? io_dataInput_122 : io_dataInput_123; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_61 = selectNodeOutputs_123 ? dataNodeOutputs_123 : dataNodeOutputs_124; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_125 = io_selectInput_124 | io_selectInput_125; // @[GameUtilities.scala 86:54]
  wire [5:0] dataNodeOutputs_125 = io_selectInput_124 ? io_dataInput_124 : io_dataInput_125; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_126 = io_selectInput_126 ? io_dataInput_126 : io_dataInput_127; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_62 = selectNodeOutputs_125 ? dataNodeOutputs_125 : dataNodeOutputs_126; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_30 = selectNodeOutputs_61 ? dataNodeOutputs_61 : dataNodeOutputs_62; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_14 = selectNodeOutputs_29 ? dataNodeOutputs_29 : dataNodeOutputs_30; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_6 = selectNodeOutputs_13 ? dataNodeOutputs_13 : dataNodeOutputs_14; // @[GameUtilities.scala 85:34]
  wire [5:0] dataNodeOutputs_2 = selectNodeOutputs_5 ? dataNodeOutputs_5 : dataNodeOutputs_6; // @[GameUtilities.scala 85:34]
  wire  selectNodeOutputs_126 = io_selectInput_126 | io_selectInput_127; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_62 = selectNodeOutputs_125 | selectNodeOutputs_126; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_30 = selectNodeOutputs_61 | selectNodeOutputs_62; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_14 = selectNodeOutputs_29 | selectNodeOutputs_30; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_6 = selectNodeOutputs_13 | selectNodeOutputs_14; // @[GameUtilities.scala 86:54]
  wire  selectNodeOutputs_2 = selectNodeOutputs_5 | selectNodeOutputs_6; // @[GameUtilities.scala 86:54]
  assign io_dataOutput = selectNodeOutputs_1 ? dataNodeOutputs_1 : dataNodeOutputs_2; // @[GameUtilities.scala 72:17]
  assign io_selectOutput = selectNodeOutputs_1 | selectNodeOutputs_2; // @[GameUtilities.scala 73:19]
endmodule
module GraphicEngineVGA(
  input         clock,
  input         reset,
  input  [10:0] io_spriteXPosition_0,
  input  [10:0] io_spriteXPosition_1,
  input  [10:0] io_spriteXPosition_2,
  input  [10:0] io_spriteXPosition_3,
  input  [10:0] io_spriteXPosition_4,
  input  [10:0] io_spriteXPosition_5,
  input  [10:0] io_spriteXPosition_6,
  input  [10:0] io_spriteXPosition_7,
  input  [10:0] io_spriteXPosition_8,
  input  [10:0] io_spriteXPosition_9,
  input  [10:0] io_spriteXPosition_10,
  input  [10:0] io_spriteXPosition_11,
  input  [10:0] io_spriteXPosition_12,
  input  [10:0] io_spriteXPosition_13,
  input  [10:0] io_spriteXPosition_14,
  input  [10:0] io_spriteXPosition_15,
  input  [10:0] io_spriteXPosition_16,
  input  [10:0] io_spriteXPosition_17,
  input  [10:0] io_spriteXPosition_18,
  input  [10:0] io_spriteXPosition_19,
  input  [10:0] io_spriteXPosition_20,
  input  [10:0] io_spriteXPosition_21,
  input  [10:0] io_spriteXPosition_22,
  input  [10:0] io_spriteXPosition_23,
  input  [10:0] io_spriteXPosition_24,
  input  [10:0] io_spriteXPosition_25,
  input  [10:0] io_spriteXPosition_26,
  input  [10:0] io_spriteXPosition_27,
  input  [10:0] io_spriteXPosition_28,
  input  [10:0] io_spriteXPosition_29,
  input  [10:0] io_spriteXPosition_30,
  input  [10:0] io_spriteXPosition_31,
  input  [10:0] io_spriteXPosition_32,
  input  [10:0] io_spriteXPosition_33,
  input  [10:0] io_spriteXPosition_41,
  input  [10:0] io_spriteXPosition_42,
  input  [10:0] io_spriteXPosition_43,
  input  [10:0] io_spriteXPosition_44,
  input  [10:0] io_spriteXPosition_45,
  input  [10:0] io_spriteXPosition_46,
  input  [10:0] io_spriteXPosition_47,
  input  [10:0] io_spriteXPosition_48,
  input  [10:0] io_spriteXPosition_49,
  input  [10:0] io_spriteXPosition_50,
  input  [10:0] io_spriteXPosition_51,
  input  [10:0] io_spriteXPosition_122,
  input  [10:0] io_spriteXPosition_123,
  input  [10:0] io_spriteXPosition_124,
  input  [10:0] io_spriteXPosition_125,
  input  [10:0] io_spriteXPosition_126,
  input  [10:0] io_spriteXPosition_127,
  input  [9:0]  io_spriteYPosition_0,
  input  [9:0]  io_spriteYPosition_1,
  input  [9:0]  io_spriteYPosition_2,
  input  [9:0]  io_spriteYPosition_3,
  input  [9:0]  io_spriteYPosition_4,
  input  [9:0]  io_spriteYPosition_5,
  input  [9:0]  io_spriteYPosition_6,
  input  [9:0]  io_spriteYPosition_7,
  input  [9:0]  io_spriteYPosition_8,
  input  [9:0]  io_spriteYPosition_9,
  input  [9:0]  io_spriteYPosition_10,
  input  [9:0]  io_spriteYPosition_11,
  input  [9:0]  io_spriteYPosition_12,
  input  [9:0]  io_spriteYPosition_13,
  input  [9:0]  io_spriteYPosition_14,
  input  [9:0]  io_spriteYPosition_15,
  input  [9:0]  io_spriteYPosition_16,
  input  [9:0]  io_spriteYPosition_17,
  input  [9:0]  io_spriteYPosition_18,
  input  [9:0]  io_spriteYPosition_19,
  input  [9:0]  io_spriteYPosition_20,
  input  [9:0]  io_spriteYPosition_21,
  input  [9:0]  io_spriteYPosition_22,
  input  [9:0]  io_spriteYPosition_23,
  input  [9:0]  io_spriteYPosition_24,
  input  [9:0]  io_spriteYPosition_25,
  input  [9:0]  io_spriteYPosition_26,
  input  [9:0]  io_spriteYPosition_27,
  input  [9:0]  io_spriteYPosition_28,
  input  [9:0]  io_spriteYPosition_29,
  input  [9:0]  io_spriteYPosition_30,
  input  [9:0]  io_spriteYPosition_31,
  input  [9:0]  io_spriteYPosition_32,
  input  [9:0]  io_spriteYPosition_33,
  input  [9:0]  io_spriteYPosition_41,
  input  [9:0]  io_spriteYPosition_42,
  input  [9:0]  io_spriteYPosition_43,
  input  [9:0]  io_spriteYPosition_122,
  input  [9:0]  io_spriteYPosition_123,
  input  [9:0]  io_spriteYPosition_124,
  input  [9:0]  io_spriteYPosition_125,
  input  [9:0]  io_spriteYPosition_126,
  input  [9:0]  io_spriteYPosition_127,
  input         io_spriteVisible_0,
  input         io_spriteVisible_1,
  input         io_spriteVisible_2,
  input         io_spriteVisible_3,
  input         io_spriteVisible_4,
  input         io_spriteVisible_5,
  input         io_spriteVisible_6,
  input         io_spriteVisible_7,
  input         io_spriteVisible_8,
  input         io_spriteVisible_9,
  input         io_spriteVisible_10,
  input         io_spriteVisible_11,
  input         io_spriteVisible_12,
  input         io_spriteVisible_13,
  input         io_spriteVisible_14,
  input         io_spriteVisible_15,
  input         io_spriteVisible_16,
  input         io_spriteVisible_17,
  input         io_spriteVisible_18,
  input         io_spriteVisible_19,
  input         io_spriteVisible_20,
  input         io_spriteVisible_21,
  input         io_spriteVisible_22,
  input         io_spriteVisible_23,
  input         io_spriteVisible_24,
  input         io_spriteVisible_25,
  input         io_spriteVisible_26,
  input         io_spriteVisible_27,
  input         io_spriteVisible_28,
  input         io_spriteVisible_29,
  input         io_spriteVisible_30,
  input         io_spriteVisible_31,
  input         io_spriteVisible_32,
  input         io_spriteVisible_33,
  input         io_spriteVisible_41,
  input         io_spriteVisible_42,
  input         io_spriteVisible_43,
  input         io_spriteVisible_44,
  input         io_spriteVisible_45,
  input         io_spriteVisible_46,
  input         io_spriteVisible_47,
  input         io_spriteVisible_48,
  input         io_spriteVisible_49,
  input         io_spriteVisible_50,
  input         io_spriteVisible_51,
  input         io_spriteVisible_55,
  input         io_spriteVisible_56,
  input         io_spriteVisible_57,
  input         io_spriteVisible_61,
  input         io_spriteVisible_62,
  input         io_spriteVisible_63,
  input         io_spriteVisible_64,
  input         io_spriteVisible_65,
  input         io_spriteVisible_66,
  input         io_spriteVisible_70,
  input         io_spriteVisible_71,
  input         io_spriteVisible_72,
  input         io_spriteFlipVertical_122,
  input         io_spriteFlipVertical_123,
  input         io_spriteFlipVertical_124,
  input         io_spriteFlipVertical_125,
  input         io_spriteFlipVertical_126,
  input         io_spriteFlipVertical_127,
  input  [9:0]  io_viewBoxX_0,
  input  [4:0]  io_backBufferWriteData,
  input  [10:0] io_backBufferWriteAddress,
  input         io_backBufferWriteEnable,
  output        io_newFrame,
  input         io_frameUpdateDone,
  output        io_missingFrameError,
  output        io_backBufferWriteError,
  output        io_viewBoxOutOfRangeError,
  output [3:0]  io_vgaRed,
  output [3:0]  io_vgaBlue,
  output [3:0]  io_vgaGreen,
  output        io_Hsync,
  output        io_Vsync
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
`endif // RANDOMIZE_REG_INIT
  wire  backTileMemories_0_0_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_0_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_0_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_1_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_1_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_1_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_2_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_2_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_2_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_3_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_3_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_3_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_4_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_4_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_4_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_5_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_5_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_5_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_6_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_6_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_6_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_7_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_7_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_7_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_8_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_8_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_8_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_9_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_9_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_9_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_10_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_10_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_10_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_11_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_11_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_11_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_12_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_12_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_12_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_13_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_13_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_13_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_14_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_14_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_14_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_15_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_15_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_15_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_16_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_16_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_16_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_17_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_17_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_17_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_18_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_18_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_18_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_19_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_19_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_19_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_20_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_20_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_20_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_21_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_21_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_21_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_22_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_22_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_22_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_23_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_23_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_23_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_24_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_24_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_24_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_25_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_25_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_25_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_26_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_26_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_26_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_27_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_27_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_27_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_28_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_28_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_28_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_29_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_29_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_29_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_30_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_30_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_30_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_0_31_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_0_31_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_0_31_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_0_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_0_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_0_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_1_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_1_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_1_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_2_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_2_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_2_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_3_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_3_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_3_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_4_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_4_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_4_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_5_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_5_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_5_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_6_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_6_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_6_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_7_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_7_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_7_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_8_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_8_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_8_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_9_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_9_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_9_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_10_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_10_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_10_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_11_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_11_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_11_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_12_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_12_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_12_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_13_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_13_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_13_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_14_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_14_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_14_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_15_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_15_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_15_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_16_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_16_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_16_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_17_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_17_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_17_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_18_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_18_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_18_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_19_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_19_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_19_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_20_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_20_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_20_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_21_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_21_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_21_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_22_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_22_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_22_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_23_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_23_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_23_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_24_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_24_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_24_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_25_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_25_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_25_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_26_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_26_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_26_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_27_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_27_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_27_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_28_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_28_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_28_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_29_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_29_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_29_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_30_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_30_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_30_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backTileMemories_1_31_clock; // @[GraphicEngineVGA.scala 162:34]
  wire [9:0] backTileMemories_1_31_io_address; // @[GraphicEngineVGA.scala 162:34]
  wire [6:0] backTileMemories_1_31_io_dataRead; // @[GraphicEngineVGA.scala 162:34]
  wire  backBufferMemories_0_clock; // @[GraphicEngineVGA.scala 186:34]
  wire [10:0] backBufferMemories_0_io_address; // @[GraphicEngineVGA.scala 186:34]
  wire [4:0] backBufferMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 186:34]
  wire  backBufferMemories_0_io_writeEnable; // @[GraphicEngineVGA.scala 186:34]
  wire [4:0] backBufferMemories_0_io_dataWrite; // @[GraphicEngineVGA.scala 186:34]
  wire  backBufferMemories_1_clock; // @[GraphicEngineVGA.scala 186:34]
  wire [10:0] backBufferMemories_1_io_address; // @[GraphicEngineVGA.scala 186:34]
  wire [4:0] backBufferMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 186:34]
  wire  backBufferMemories_1_io_writeEnable; // @[GraphicEngineVGA.scala 186:34]
  wire [4:0] backBufferMemories_1_io_dataWrite; // @[GraphicEngineVGA.scala 186:34]
  wire  backBufferShadowMemories_0_clock; // @[GraphicEngineVGA.scala 191:40]
  wire [10:0] backBufferShadowMemories_0_io_address; // @[GraphicEngineVGA.scala 191:40]
  wire [4:0] backBufferShadowMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 191:40]
  wire  backBufferShadowMemories_0_io_writeEnable; // @[GraphicEngineVGA.scala 191:40]
  wire [4:0] backBufferShadowMemories_0_io_dataWrite; // @[GraphicEngineVGA.scala 191:40]
  wire  backBufferShadowMemories_1_clock; // @[GraphicEngineVGA.scala 191:40]
  wire [10:0] backBufferShadowMemories_1_io_address; // @[GraphicEngineVGA.scala 191:40]
  wire [4:0] backBufferShadowMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 191:40]
  wire  backBufferShadowMemories_1_io_writeEnable; // @[GraphicEngineVGA.scala 191:40]
  wire [4:0] backBufferShadowMemories_1_io_dataWrite; // @[GraphicEngineVGA.scala 191:40]
  wire  backBufferRestoreMemories_0_clock; // @[GraphicEngineVGA.scala 197:41]
  wire [10:0] backBufferRestoreMemories_0_io_address; // @[GraphicEngineVGA.scala 197:41]
  wire [4:0] backBufferRestoreMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 197:41]
  wire  backBufferRestoreMemories_1_clock; // @[GraphicEngineVGA.scala 197:41]
  wire [10:0] backBufferRestoreMemories_1_io_address; // @[GraphicEngineVGA.scala 197:41]
  wire [4:0] backBufferRestoreMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 197:41]
  wire  spriteMemories_0_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_0_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_1_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_1_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_2_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_2_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_2_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_3_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_3_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_3_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_4_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_4_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_4_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_5_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_5_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_5_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_6_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_6_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_6_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_7_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_7_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_7_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_8_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_8_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_8_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_9_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_9_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_9_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_10_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_10_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_10_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_11_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_11_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_11_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_12_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_12_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_12_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_13_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_13_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_13_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_14_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_14_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_14_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_15_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_15_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_15_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_16_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_16_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_16_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_17_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_17_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_17_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_18_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_18_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_18_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_19_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_19_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_19_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_20_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_20_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_20_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_21_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_21_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_21_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_22_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_22_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_22_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_23_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_23_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_23_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_24_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_24_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_24_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_25_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_25_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_25_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_26_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_26_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_26_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_27_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_27_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_27_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_28_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_28_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_28_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_29_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_29_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_29_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_30_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_30_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_30_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_31_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_31_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_31_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_32_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_32_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_32_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_33_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_33_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_33_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_34_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_34_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_34_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_35_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_35_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_35_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_36_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_36_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_36_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_37_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_37_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_37_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_38_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_38_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_38_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_39_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_39_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_39_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_40_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_40_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_40_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_41_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_41_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_41_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_42_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_42_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_42_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_43_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_43_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_43_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_44_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_44_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_44_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_45_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_45_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_45_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_46_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_46_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_46_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_47_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_47_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_47_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_48_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_48_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_48_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_49_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_49_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_49_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_50_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_50_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_50_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_51_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_51_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_51_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_52_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_52_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_52_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_53_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_53_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_53_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_54_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_54_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_54_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_55_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_55_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_55_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_56_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_56_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_56_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_57_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_57_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_57_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_58_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_58_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_58_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_59_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_59_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_59_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_60_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_60_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_60_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_61_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_61_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_61_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_62_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_62_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_62_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_63_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_63_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_63_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_64_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_64_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_64_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_65_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_65_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_65_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_66_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_66_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_66_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_67_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_67_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_67_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_68_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_68_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_68_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_69_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_69_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_69_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_70_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_70_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_70_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_71_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_71_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_71_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_72_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_72_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_72_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_73_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_73_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_73_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_74_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_74_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_74_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_75_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_75_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_75_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_76_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_76_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_76_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_77_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_77_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_77_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_78_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_78_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_78_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_79_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_79_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_79_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_80_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_80_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_80_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_81_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_81_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_81_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_82_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_82_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_82_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_83_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_83_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_83_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_84_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_84_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_84_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_85_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_85_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_85_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_86_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_86_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_86_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_87_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_87_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_87_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_88_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_88_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_88_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_89_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_89_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_89_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_90_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_90_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_90_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_91_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_91_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_91_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_92_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_92_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_92_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_93_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_93_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_93_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_94_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_94_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_94_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_95_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_95_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_95_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_96_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_96_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_96_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_97_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_97_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_97_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_98_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_98_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_98_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_99_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_99_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_99_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_100_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_100_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_100_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_101_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_101_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_101_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_102_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_102_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_102_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_103_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_103_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_103_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_104_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_104_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_104_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_105_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_105_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_105_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_106_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_106_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_106_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_107_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_107_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_107_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_108_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_108_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_108_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_109_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_109_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_109_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_110_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_110_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_110_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_111_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_111_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_111_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_112_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_112_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_112_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_113_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_113_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_113_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_114_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_114_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_114_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_115_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_115_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_115_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_116_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_116_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_116_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_117_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_117_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_117_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_118_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_118_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_118_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_119_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_119_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_119_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_120_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_120_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_120_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_121_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_121_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_121_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_122_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_122_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_122_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_123_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_123_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_123_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_124_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_124_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_124_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_125_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_125_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_125_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_126_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_126_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_126_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire  spriteMemories_127_clock; // @[GraphicEngineVGA.scala 273:30]
  wire [9:0] spriteMemories_127_io_address; // @[GraphicEngineVGA.scala 273:30]
  wire [6:0] spriteMemories_127_io_dataRead; // @[GraphicEngineVGA.scala 273:30]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_0; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_1; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_2; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_3; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_4; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_5; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_6; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_7; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_8; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_9; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_10; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_11; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_12; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_13; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_14; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_15; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_16; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_17; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_18; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_19; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_20; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_21; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_22; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_23; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_24; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_25; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_26; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_27; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_28; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_29; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_30; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_31; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_32; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_33; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_34; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_35; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_36; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_37; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_38; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_39; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_40; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_41; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_42; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_43; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_44; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_45; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_46; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_47; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_48; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_49; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_50; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_51; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_52; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_53; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_54; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_55; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_56; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_57; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_58; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_59; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_60; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_61; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_62; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_63; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_64; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_65; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_66; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_67; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_68; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_69; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_70; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_71; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_72; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_73; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_74; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_75; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_76; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_77; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_78; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_79; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_80; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_81; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_82; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_83; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_84; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_85; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_86; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_87; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_88; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_89; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_90; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_91; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_92; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_93; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_94; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_95; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_96; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_97; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_98; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_99; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_100; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_101; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_102; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_103; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_104; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_105; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_106; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_107; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_108; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_109; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_110; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_111; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_112; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_113; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_114; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_115; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_116; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_117; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_118; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_119; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_120; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_121; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_122; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_123; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_124; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_125; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_126; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataInput_127; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_0; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_1; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_2; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_3; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_4; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_5; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_6; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_7; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_8; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_9; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_10; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_11; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_12; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_13; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_14; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_15; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_16; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_17; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_18; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_19; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_20; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_21; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_22; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_23; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_24; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_25; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_26; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_27; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_28; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_29; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_30; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_31; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_32; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_33; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_34; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_35; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_36; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_37; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_38; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_39; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_40; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_41; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_42; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_43; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_44; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_45; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_46; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_47; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_48; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_49; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_50; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_51; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_52; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_53; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_54; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_55; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_56; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_57; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_58; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_59; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_60; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_61; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_62; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_63; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_64; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_65; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_66; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_67; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_68; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_69; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_70; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_71; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_72; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_73; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_74; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_75; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_76; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_77; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_78; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_79; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_80; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_81; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_82; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_83; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_84; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_85; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_86; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_87; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_88; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_89; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_90; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_91; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_92; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_93; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_94; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_95; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_96; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_97; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_98; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_99; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_100; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_101; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_102; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_103; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_104; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_105; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_106; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_107; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_108; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_109; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_110; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_111; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_112; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_113; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_114; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_115; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_116; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_117; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_118; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_119; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_120; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_121; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_122; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_123; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_124; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_125; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_126; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectInput_127; // @[GraphicEngineVGA.scala 306:44]
  wire [5:0] multiHotPriortyReductionTree_io_dataOutput; // @[GraphicEngineVGA.scala 306:44]
  wire  multiHotPriortyReductionTree_io_selectOutput; // @[GraphicEngineVGA.scala 306:44]
  reg [1:0] ScaleCounterReg; // @[GraphicEngineVGA.scala 63:32]
  reg [9:0] CounterXReg; // @[GraphicEngineVGA.scala 64:28]
  reg [9:0] CounterYReg; // @[GraphicEngineVGA.scala 65:28]
  wire  _T = ScaleCounterReg == 2'h3; // @[GraphicEngineVGA.scala 70:26]
  wire  _T_1 = CounterXReg == 10'h31f; // @[GraphicEngineVGA.scala 72:24]
  wire  _T_2 = CounterYReg == 10'h20c; // @[GraphicEngineVGA.scala 74:26]
  wire [9:0] _T_4 = CounterYReg + 10'h1; // @[GraphicEngineVGA.scala 78:38]
  wire [9:0] _T_6 = CounterXReg + 10'h1; // @[GraphicEngineVGA.scala 81:36]
  wire  _GEN_4 = _T_1 & _T_2; // @[GraphicEngineVGA.scala 72:129]
  wire [1:0] _T_8 = ScaleCounterReg + 2'h1; // @[GraphicEngineVGA.scala 84:42]
  wire  _GEN_8 = _T & _GEN_4; // @[GraphicEngineVGA.scala 70:52]
  reg [11:0] backMemoryRestoreCounter; // @[GraphicEngineVGA.scala 220:41]
  wire  restoreEnabled = backMemoryRestoreCounter < 12'h800; // @[GraphicEngineVGA.scala 223:33]
  wire  run = restoreEnabled ? 1'h0 : 1'h1; // @[GraphicEngineVGA.scala 223:70]
  wire  _T_9 = CounterXReg >= 10'h290; // @[GraphicEngineVGA.scala 88:28]
  wire  _T_10 = CounterXReg < 10'h2f0; // @[GraphicEngineVGA.scala 88:95]
  wire  Hsync = _T_9 & _T_10; // @[GraphicEngineVGA.scala 88:79]
  wire  _T_11 = CounterYReg >= 10'h1ea; // @[GraphicEngineVGA.scala 89:28]
  wire  _T_12 = CounterYReg < 10'h1ec; // @[GraphicEngineVGA.scala 89:95]
  wire  Vsync = _T_11 & _T_12; // @[GraphicEngineVGA.scala 89:79]
  reg  _T_14_0; // @[GameUtilities.scala 21:24]
  reg  _T_14_1; // @[GameUtilities.scala 21:24]
  reg  _T_14_2; // @[GameUtilities.scala 21:24]
  reg  _T_14_3; // @[GameUtilities.scala 21:24]
  reg  _T_16_0; // @[GameUtilities.scala 21:24]
  reg  _T_16_1; // @[GameUtilities.scala 21:24]
  reg  _T_16_2; // @[GameUtilities.scala 21:24]
  reg  _T_16_3; // @[GameUtilities.scala 21:24]
  wire  _T_17 = CounterXReg < 10'h280; // @[GraphicEngineVGA.scala 93:36]
  wire  _T_18 = CounterYReg < 10'h1e0; // @[GraphicEngineVGA.scala 93:76]
  reg [20:0] frameClockCount; // @[GraphicEngineVGA.scala 100:32]
  wire  _T_19 = frameClockCount == 21'h19a27f; // @[GraphicEngineVGA.scala 101:42]
  wire [20:0] _T_21 = frameClockCount + 21'h1; // @[GraphicEngineVGA.scala 101:92]
  wire  preDisplayArea = frameClockCount >= 21'h199a1b; // @[GraphicEngineVGA.scala 102:40]
  reg [10:0] spriteXPositionReg_0; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_1; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_2; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_3; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_4; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_5; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_6; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_7; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_8; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_9; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_10; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_11; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_12; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_13; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_14; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_15; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_16; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_17; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_18; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_19; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_20; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_21; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_22; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_23; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_24; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_25; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_26; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_27; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_28; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_29; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_30; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_31; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_32; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_33; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_34; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_35; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_36; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_37; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_38; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_39; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_40; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_41; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_42; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_43; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_44; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_45; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_46; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_47; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_48; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_49; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_50; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_51; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_52; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_53; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_54; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_55; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_56; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_57; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_58; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_59; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_60; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_61; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_62; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_63; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_64; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_65; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_66; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_67; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_68; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_69; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_70; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_71; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_72; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_73; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_74; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_75; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_76; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_77; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_78; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_79; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_80; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_81; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_82; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_83; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_84; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_85; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_86; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_87; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_88; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_89; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_90; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_91; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_92; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_93; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_94; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_95; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_96; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_97; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_98; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_99; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_100; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_101; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_102; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_103; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_104; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_105; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_106; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_107; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_108; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_109; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_110; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_111; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_112; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_113; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_114; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_115; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_116; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_117; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_118; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_119; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_120; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_121; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_122; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_123; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_124; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_125; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_126; // @[Reg.scala 27:20]
  reg [10:0] spriteXPositionReg_127; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_0; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_1; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_2; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_3; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_4; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_5; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_6; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_7; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_8; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_9; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_10; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_11; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_12; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_13; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_14; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_15; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_16; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_17; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_18; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_19; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_20; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_21; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_22; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_23; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_24; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_25; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_26; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_27; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_28; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_29; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_30; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_31; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_32; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_33; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_34; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_35; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_36; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_37; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_38; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_39; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_40; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_41; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_42; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_43; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_44; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_45; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_46; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_47; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_48; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_49; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_50; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_51; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_52; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_53; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_54; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_55; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_56; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_57; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_58; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_59; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_60; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_61; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_62; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_63; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_70; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_71; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_72; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_73; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_74; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_75; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_76; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_77; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_78; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_79; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_80; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_81; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_82; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_83; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_84; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_85; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_86; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_87; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_88; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_89; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_90; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_91; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_92; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_93; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_94; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_95; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_96; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_97; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_98; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_99; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_100; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_101; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_102; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_103; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_104; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_105; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_106; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_107; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_108; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_109; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_110; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_111; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_112; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_113; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_114; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_115; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_116; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_117; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_118; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_119; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_120; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_121; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_122; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_123; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_124; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_125; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_126; // @[Reg.scala 27:20]
  reg [9:0] spriteYPositionReg_127; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_0; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_1; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_2; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_3; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_4; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_5; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_6; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_7; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_8; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_9; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_10; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_11; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_12; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_13; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_14; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_15; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_16; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_17; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_18; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_19; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_20; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_21; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_22; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_23; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_24; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_25; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_26; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_27; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_28; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_29; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_30; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_31; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_32; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_33; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_41; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_42; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_43; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_44; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_45; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_46; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_47; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_48; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_49; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_50; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_51; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_55; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_56; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_57; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_61; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_62; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_63; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_64; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_65; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_66; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_70; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_71; // @[Reg.scala 27:20]
  reg  spriteVisibleReg_72; // @[Reg.scala 27:20]
  wire  _GEN_269 = io_newFrame ? io_spriteVisible_0 : spriteVisibleReg_0; // @[Reg.scala 28:19]
  wire  _GEN_270 = io_newFrame ? io_spriteVisible_1 : spriteVisibleReg_1; // @[Reg.scala 28:19]
  wire  _GEN_271 = io_newFrame ? io_spriteVisible_2 : spriteVisibleReg_2; // @[Reg.scala 28:19]
  wire  _GEN_272 = io_newFrame ? io_spriteVisible_3 : spriteVisibleReg_3; // @[Reg.scala 28:19]
  wire  _GEN_273 = io_newFrame ? io_spriteVisible_4 : spriteVisibleReg_4; // @[Reg.scala 28:19]
  wire  _GEN_274 = io_newFrame ? io_spriteVisible_5 : spriteVisibleReg_5; // @[Reg.scala 28:19]
  wire  _GEN_275 = io_newFrame ? io_spriteVisible_6 : spriteVisibleReg_6; // @[Reg.scala 28:19]
  wire  _GEN_276 = io_newFrame ? io_spriteVisible_7 : spriteVisibleReg_7; // @[Reg.scala 28:19]
  wire  _GEN_277 = io_newFrame ? io_spriteVisible_8 : spriteVisibleReg_8; // @[Reg.scala 28:19]
  wire  _GEN_278 = io_newFrame ? io_spriteVisible_9 : spriteVisibleReg_9; // @[Reg.scala 28:19]
  wire  _GEN_279 = io_newFrame ? io_spriteVisible_10 : spriteVisibleReg_10; // @[Reg.scala 28:19]
  wire  _GEN_280 = io_newFrame ? io_spriteVisible_11 : spriteVisibleReg_11; // @[Reg.scala 28:19]
  wire  _GEN_281 = io_newFrame ? io_spriteVisible_12 : spriteVisibleReg_12; // @[Reg.scala 28:19]
  wire  _GEN_282 = io_newFrame ? io_spriteVisible_13 : spriteVisibleReg_13; // @[Reg.scala 28:19]
  wire  _GEN_283 = io_newFrame ? io_spriteVisible_14 : spriteVisibleReg_14; // @[Reg.scala 28:19]
  wire  _GEN_284 = io_newFrame ? io_spriteVisible_15 : spriteVisibleReg_15; // @[Reg.scala 28:19]
  wire  _GEN_285 = io_newFrame ? io_spriteVisible_16 : spriteVisibleReg_16; // @[Reg.scala 28:19]
  wire  _GEN_286 = io_newFrame ? io_spriteVisible_17 : spriteVisibleReg_17; // @[Reg.scala 28:19]
  wire  _GEN_287 = io_newFrame ? io_spriteVisible_18 : spriteVisibleReg_18; // @[Reg.scala 28:19]
  wire  _GEN_288 = io_newFrame ? io_spriteVisible_19 : spriteVisibleReg_19; // @[Reg.scala 28:19]
  wire  _GEN_289 = io_newFrame ? io_spriteVisible_20 : spriteVisibleReg_20; // @[Reg.scala 28:19]
  wire  _GEN_290 = io_newFrame ? io_spriteVisible_21 : spriteVisibleReg_21; // @[Reg.scala 28:19]
  wire  _GEN_291 = io_newFrame ? io_spriteVisible_22 : spriteVisibleReg_22; // @[Reg.scala 28:19]
  wire  _GEN_292 = io_newFrame ? io_spriteVisible_23 : spriteVisibleReg_23; // @[Reg.scala 28:19]
  wire  _GEN_293 = io_newFrame ? io_spriteVisible_24 : spriteVisibleReg_24; // @[Reg.scala 28:19]
  wire  _GEN_294 = io_newFrame ? io_spriteVisible_25 : spriteVisibleReg_25; // @[Reg.scala 28:19]
  wire  _GEN_295 = io_newFrame ? io_spriteVisible_26 : spriteVisibleReg_26; // @[Reg.scala 28:19]
  wire  _GEN_296 = io_newFrame ? io_spriteVisible_27 : spriteVisibleReg_27; // @[Reg.scala 28:19]
  wire  _GEN_297 = io_newFrame ? io_spriteVisible_28 : spriteVisibleReg_28; // @[Reg.scala 28:19]
  wire  _GEN_298 = io_newFrame ? io_spriteVisible_29 : spriteVisibleReg_29; // @[Reg.scala 28:19]
  wire  _GEN_299 = io_newFrame ? io_spriteVisible_30 : spriteVisibleReg_30; // @[Reg.scala 28:19]
  wire  _GEN_300 = io_newFrame ? io_spriteVisible_31 : spriteVisibleReg_31; // @[Reg.scala 28:19]
  wire  _GEN_301 = io_newFrame ? io_spriteVisible_32 : spriteVisibleReg_32; // @[Reg.scala 28:19]
  wire  _GEN_302 = io_newFrame ? io_spriteVisible_33 : spriteVisibleReg_33; // @[Reg.scala 28:19]
  wire  _GEN_310 = io_newFrame ? io_spriteVisible_41 : spriteVisibleReg_41; // @[Reg.scala 28:19]
  wire  _GEN_311 = io_newFrame ? io_spriteVisible_42 : spriteVisibleReg_42; // @[Reg.scala 28:19]
  wire  _GEN_312 = io_newFrame ? io_spriteVisible_43 : spriteVisibleReg_43; // @[Reg.scala 28:19]
  wire  _GEN_313 = io_newFrame ? io_spriteVisible_44 : spriteVisibleReg_44; // @[Reg.scala 28:19]
  wire  _GEN_314 = io_newFrame ? io_spriteVisible_45 : spriteVisibleReg_45; // @[Reg.scala 28:19]
  wire  _GEN_315 = io_newFrame ? io_spriteVisible_46 : spriteVisibleReg_46; // @[Reg.scala 28:19]
  wire  _GEN_316 = io_newFrame ? io_spriteVisible_47 : spriteVisibleReg_47; // @[Reg.scala 28:19]
  wire  _GEN_317 = io_newFrame ? io_spriteVisible_48 : spriteVisibleReg_48; // @[Reg.scala 28:19]
  wire  _GEN_318 = io_newFrame ? io_spriteVisible_49 : spriteVisibleReg_49; // @[Reg.scala 28:19]
  wire  _GEN_319 = io_newFrame ? io_spriteVisible_50 : spriteVisibleReg_50; // @[Reg.scala 28:19]
  wire  _GEN_320 = io_newFrame ? io_spriteVisible_51 : spriteVisibleReg_51; // @[Reg.scala 28:19]
  wire  _GEN_324 = io_newFrame ? io_spriteVisible_55 : spriteVisibleReg_55; // @[Reg.scala 28:19]
  wire  _GEN_325 = io_newFrame ? io_spriteVisible_56 : spriteVisibleReg_56; // @[Reg.scala 28:19]
  wire  _GEN_326 = io_newFrame ? io_spriteVisible_57 : spriteVisibleReg_57; // @[Reg.scala 28:19]
  wire  _GEN_330 = io_newFrame ? io_spriteVisible_61 : spriteVisibleReg_61; // @[Reg.scala 28:19]
  wire  _GEN_331 = io_newFrame ? io_spriteVisible_62 : spriteVisibleReg_62; // @[Reg.scala 28:19]
  wire  _GEN_332 = io_newFrame ? io_spriteVisible_63 : spriteVisibleReg_63; // @[Reg.scala 28:19]
  wire  _GEN_333 = io_newFrame ? io_spriteVisible_64 : spriteVisibleReg_64; // @[Reg.scala 28:19]
  wire  _GEN_334 = io_newFrame ? io_spriteVisible_65 : spriteVisibleReg_65; // @[Reg.scala 28:19]
  wire  _GEN_335 = io_newFrame ? io_spriteVisible_66 : spriteVisibleReg_66; // @[Reg.scala 28:19]
  wire  _GEN_339 = io_newFrame ? io_spriteVisible_70 : spriteVisibleReg_70; // @[Reg.scala 28:19]
  wire  _GEN_340 = io_newFrame ? io_spriteVisible_71 : spriteVisibleReg_71; // @[Reg.scala 28:19]
  wire  _GEN_341 = io_newFrame ? io_spriteVisible_72 : spriteVisibleReg_72; // @[Reg.scala 28:19]
  reg  spriteFlipVerticalReg_122; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_123; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_124; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_125; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_126; // @[Reg.scala 27:20]
  reg  spriteFlipVerticalReg_127; // @[Reg.scala 27:20]
  reg [9:0] viewBoxXReg_0; // @[Reg.scala 27:20]
  reg  missingFrameErrorReg; // @[GraphicEngineVGA.scala 122:37]
  reg  backBufferWriteErrorReg; // @[GraphicEngineVGA.scala 123:40]
  reg  viewBoxOutOfRangeErrorReg; // @[GraphicEngineVGA.scala 124:42]
  wire  _T_28 = viewBoxXReg_0 >= 10'h280; // @[GraphicEngineVGA.scala 136:45]
  wire [9:0] viewBoxXClipped_0 = _T_28 ? 10'h280 : viewBoxXReg_0; // @[GraphicEngineVGA.scala 136:29]
  wire [10:0] pixelXBack_0 = CounterXReg + viewBoxXClipped_0; // @[GraphicEngineVGA.scala 138:29]
  wire [10:0] pixelYBack_0 = {{1'd0}, CounterYReg}; // @[GraphicEngineVGA.scala 139:29]
  wire [10:0] pixelXBack_1 = {{1'd0}, CounterXReg}; // @[GraphicEngineVGA.scala 138:29]
  wire  _T_40 = viewBoxXReg_0 > 10'h280; // @[GraphicEngineVGA.scala 142:23]
  wire  _GEN_657 = _T_40 | viewBoxOutOfRangeErrorReg; // @[GraphicEngineVGA.scala 142:58]
  reg  newFrameStikyReg; // @[GraphicEngineVGA.scala 149:33]
  wire  _GEN_658 = io_newFrame | newFrameStikyReg; // @[GraphicEngineVGA.scala 150:21]
  reg  _T_43; // @[GraphicEngineVGA.scala 153:16]
  wire  _T_44 = newFrameStikyReg & io_newFrame; // @[GraphicEngineVGA.scala 156:26]
  wire  _GEN_660 = _T_44 | missingFrameErrorReg; // @[GraphicEngineVGA.scala 156:41]
  wire [5:0] _GEN_990 = {{1'd0}, pixelYBack_0[4:0]}; // @[GraphicEngineVGA.scala 175:82]
  wire [10:0] _T_47 = 6'h20 * _GEN_990; // @[GraphicEngineVGA.scala 175:82]
  wire [10:0] _GEN_991 = {{6'd0}, pixelXBack_0[4:0]}; // @[GraphicEngineVGA.scala 175:69]
  wire [11:0] _T_48 = _GEN_991 + _T_47; // @[GraphicEngineVGA.scala 175:69]
  reg [6:0] backTileMemoryDataRead_0_0; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_1; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_2; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_3; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_4; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_5; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_6; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_7; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_8; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_9; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_10; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_11; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_12; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_13; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_14; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_15; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_16; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_17; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_18; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_19; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_20; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_21; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_22; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_23; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_24; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_25; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_26; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_27; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_28; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_29; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_30; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_0_31; // @[GraphicEngineVGA.scala 177:44]
  wire [10:0] _GEN_1055 = {{6'd0}, pixelXBack_1[4:0]}; // @[GraphicEngineVGA.scala 175:69]
  wire [11:0] _T_208 = _GEN_1055 + _T_47; // @[GraphicEngineVGA.scala 175:69]
  reg [6:0] backTileMemoryDataRead_1_0; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_1; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_2; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_3; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_4; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_5; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_6; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_7; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_8; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_9; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_10; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_11; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_12; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_13; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_14; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_15; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_16; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_17; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_18; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_19; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_20; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_21; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_22; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_23; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_24; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_25; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_26; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_27; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_28; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_29; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_30; // @[GraphicEngineVGA.scala 177:44]
  reg [6:0] backTileMemoryDataRead_1_31; // @[GraphicEngineVGA.scala 177:44]
  reg [11:0] backMemoryCopyCounter; // @[GraphicEngineVGA.scala 201:38]
  wire  _T_365 = backMemoryCopyCounter < 12'h800; // @[GraphicEngineVGA.scala 205:32]
  wire [11:0] _T_367 = backMemoryCopyCounter + 12'h1; // @[GraphicEngineVGA.scala 206:54]
  wire  copyEnabled = preDisplayArea & _T_365; // @[GraphicEngineVGA.scala 204:23]
  reg  copyEnabledReg; // @[GraphicEngineVGA.scala 218:31]
  wire [11:0] _T_370 = backMemoryRestoreCounter + 12'h1; // @[GraphicEngineVGA.scala 224:58]
  reg [10:0] _T_373; // @[GraphicEngineVGA.scala 240:72]
  reg [10:0] _T_375; // @[GraphicEngineVGA.scala 240:161]
  wire [10:0] _T_376 = copyEnabled ? backMemoryCopyCounter[10:0] : _T_375; // @[GraphicEngineVGA.scala 240:110]
  reg  _T_378; // @[GraphicEngineVGA.scala 242:76]
  reg  _T_379; // @[GraphicEngineVGA.scala 242:127]
  wire  _T_380 = copyEnabled ? 1'h0 : _T_379; // @[GraphicEngineVGA.scala 242:97]
  reg [4:0] _T_382; // @[GraphicEngineVGA.scala 243:116]
  reg [10:0] _T_385; // @[GraphicEngineVGA.scala 245:66]
  wire [11:0] _T_388 = 6'h28 * pixelYBack_0[10:5]; // @[GraphicEngineVGA.scala 245:139]
  wire [11:0] _GEN_1118 = {{6'd0}, pixelXBack_0[10:5]}; // @[GraphicEngineVGA.scala 245:126]
  wire [12:0] _T_389 = _GEN_1118 + _T_388; // @[GraphicEngineVGA.scala 245:126]
  wire [12:0] _T_390 = copyEnabledReg ? {{2'd0}, _T_385} : _T_389; // @[GraphicEngineVGA.scala 245:42]
  reg [10:0] _T_393; // @[GraphicEngineVGA.scala 240:72]
  reg [10:0] _T_395; // @[GraphicEngineVGA.scala 240:161]
  wire [10:0] _T_396 = copyEnabled ? backMemoryCopyCounter[10:0] : _T_395; // @[GraphicEngineVGA.scala 240:110]
  reg  _T_398; // @[GraphicEngineVGA.scala 242:76]
  reg  _T_399; // @[GraphicEngineVGA.scala 242:127]
  wire  _T_400 = copyEnabled ? 1'h0 : _T_399; // @[GraphicEngineVGA.scala 242:97]
  reg [4:0] _T_402; // @[GraphicEngineVGA.scala 243:116]
  reg [10:0] _T_405; // @[GraphicEngineVGA.scala 245:66]
  wire [11:0] _GEN_1119 = {{6'd0}, pixelXBack_1[10:5]}; // @[GraphicEngineVGA.scala 245:126]
  wire [12:0] _T_409 = _GEN_1119 + _T_388; // @[GraphicEngineVGA.scala 245:126]
  wire [12:0] _T_410 = copyEnabledReg ? {{2'd0}, _T_405} : _T_409; // @[GraphicEngineVGA.scala 245:42]
  wire  _T_411 = copyEnabled | copyEnabledReg; // @[GraphicEngineVGA.scala 252:20]
  wire  _GEN_668 = io_backBufferWriteEnable | backBufferWriteErrorReg; // @[GraphicEngineVGA.scala 253:36]
  reg [4:0] _T_412; // @[GraphicEngineVGA.scala 265:64]
  wire [6:0] _GEN_671 = 5'h1 == _T_412 ? backTileMemoryDataRead_0_1 : backTileMemoryDataRead_0_0; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_672 = 5'h2 == _T_412 ? backTileMemoryDataRead_0_2 : _GEN_671; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_673 = 5'h3 == _T_412 ? backTileMemoryDataRead_0_3 : _GEN_672; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_674 = 5'h4 == _T_412 ? backTileMemoryDataRead_0_4 : _GEN_673; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_675 = 5'h5 == _T_412 ? backTileMemoryDataRead_0_5 : _GEN_674; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_676 = 5'h6 == _T_412 ? backTileMemoryDataRead_0_6 : _GEN_675; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_677 = 5'h7 == _T_412 ? backTileMemoryDataRead_0_7 : _GEN_676; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_678 = 5'h8 == _T_412 ? backTileMemoryDataRead_0_8 : _GEN_677; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_679 = 5'h9 == _T_412 ? backTileMemoryDataRead_0_9 : _GEN_678; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_680 = 5'ha == _T_412 ? backTileMemoryDataRead_0_10 : _GEN_679; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_681 = 5'hb == _T_412 ? backTileMemoryDataRead_0_11 : _GEN_680; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_682 = 5'hc == _T_412 ? backTileMemoryDataRead_0_12 : _GEN_681; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_683 = 5'hd == _T_412 ? backTileMemoryDataRead_0_13 : _GEN_682; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_684 = 5'he == _T_412 ? backTileMemoryDataRead_0_14 : _GEN_683; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_685 = 5'hf == _T_412 ? backTileMemoryDataRead_0_15 : _GEN_684; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_686 = 5'h10 == _T_412 ? backTileMemoryDataRead_0_16 : _GEN_685; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_687 = 5'h11 == _T_412 ? backTileMemoryDataRead_0_17 : _GEN_686; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_688 = 5'h12 == _T_412 ? backTileMemoryDataRead_0_18 : _GEN_687; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_689 = 5'h13 == _T_412 ? backTileMemoryDataRead_0_19 : _GEN_688; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_690 = 5'h14 == _T_412 ? backTileMemoryDataRead_0_20 : _GEN_689; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_691 = 5'h15 == _T_412 ? backTileMemoryDataRead_0_21 : _GEN_690; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_692 = 5'h16 == _T_412 ? backTileMemoryDataRead_0_22 : _GEN_691; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_693 = 5'h17 == _T_412 ? backTileMemoryDataRead_0_23 : _GEN_692; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_694 = 5'h18 == _T_412 ? backTileMemoryDataRead_0_24 : _GEN_693; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_695 = 5'h19 == _T_412 ? backTileMemoryDataRead_0_25 : _GEN_694; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_696 = 5'h1a == _T_412 ? backTileMemoryDataRead_0_26 : _GEN_695; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_697 = 5'h1b == _T_412 ? backTileMemoryDataRead_0_27 : _GEN_696; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_698 = 5'h1c == _T_412 ? backTileMemoryDataRead_0_28 : _GEN_697; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_699 = 5'h1d == _T_412 ? backTileMemoryDataRead_0_29 : _GEN_698; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_700 = 5'h1e == _T_412 ? backTileMemoryDataRead_0_30 : _GEN_699; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] fullBackgroundColor_0 = 5'h1f == _T_412 ? backTileMemoryDataRead_0_31 : _GEN_700; // @[GraphicEngineVGA.scala 265:28]
  reg [4:0] _T_415; // @[GraphicEngineVGA.scala 265:64]
  wire [6:0] _GEN_703 = 5'h1 == _T_415 ? backTileMemoryDataRead_1_1 : backTileMemoryDataRead_1_0; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_704 = 5'h2 == _T_415 ? backTileMemoryDataRead_1_2 : _GEN_703; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_705 = 5'h3 == _T_415 ? backTileMemoryDataRead_1_3 : _GEN_704; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_706 = 5'h4 == _T_415 ? backTileMemoryDataRead_1_4 : _GEN_705; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_707 = 5'h5 == _T_415 ? backTileMemoryDataRead_1_5 : _GEN_706; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_708 = 5'h6 == _T_415 ? backTileMemoryDataRead_1_6 : _GEN_707; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_709 = 5'h7 == _T_415 ? backTileMemoryDataRead_1_7 : _GEN_708; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_710 = 5'h8 == _T_415 ? backTileMemoryDataRead_1_8 : _GEN_709; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_711 = 5'h9 == _T_415 ? backTileMemoryDataRead_1_9 : _GEN_710; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_712 = 5'ha == _T_415 ? backTileMemoryDataRead_1_10 : _GEN_711; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_713 = 5'hb == _T_415 ? backTileMemoryDataRead_1_11 : _GEN_712; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_714 = 5'hc == _T_415 ? backTileMemoryDataRead_1_12 : _GEN_713; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_715 = 5'hd == _T_415 ? backTileMemoryDataRead_1_13 : _GEN_714; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_716 = 5'he == _T_415 ? backTileMemoryDataRead_1_14 : _GEN_715; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_717 = 5'hf == _T_415 ? backTileMemoryDataRead_1_15 : _GEN_716; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_718 = 5'h10 == _T_415 ? backTileMemoryDataRead_1_16 : _GEN_717; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_719 = 5'h11 == _T_415 ? backTileMemoryDataRead_1_17 : _GEN_718; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_720 = 5'h12 == _T_415 ? backTileMemoryDataRead_1_18 : _GEN_719; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_721 = 5'h13 == _T_415 ? backTileMemoryDataRead_1_19 : _GEN_720; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_722 = 5'h14 == _T_415 ? backTileMemoryDataRead_1_20 : _GEN_721; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_723 = 5'h15 == _T_415 ? backTileMemoryDataRead_1_21 : _GEN_722; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_724 = 5'h16 == _T_415 ? backTileMemoryDataRead_1_22 : _GEN_723; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_725 = 5'h17 == _T_415 ? backTileMemoryDataRead_1_23 : _GEN_724; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_726 = 5'h18 == _T_415 ? backTileMemoryDataRead_1_24 : _GEN_725; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_727 = 5'h19 == _T_415 ? backTileMemoryDataRead_1_25 : _GEN_726; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_728 = 5'h1a == _T_415 ? backTileMemoryDataRead_1_26 : _GEN_727; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_729 = 5'h1b == _T_415 ? backTileMemoryDataRead_1_27 : _GEN_728; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_730 = 5'h1c == _T_415 ? backTileMemoryDataRead_1_28 : _GEN_729; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_731 = 5'h1d == _T_415 ? backTileMemoryDataRead_1_29 : _GEN_730; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] _GEN_732 = 5'h1e == _T_415 ? backTileMemoryDataRead_1_30 : _GEN_731; // @[GraphicEngineVGA.scala 265:28]
  wire [6:0] fullBackgroundColor_1 = 5'h1f == _T_415 ? backTileMemoryDataRead_1_31 : _GEN_732; // @[GraphicEngineVGA.scala 265:28]
  reg [5:0] pixelColorBack; // @[GraphicEngineVGA.scala 268:31]
  wire [10:0] _T_425 = {1'h0,CounterXReg}; // @[GraphicEngineVGA.scala 281:47]
  wire [11:0] inSpriteX_0 = $signed(_T_425) - $signed(spriteXPositionReg_0); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _T_431 = {1'h0,CounterYReg}; // @[GraphicEngineVGA.scala 287:47]
  wire [10:0] _GEN_1120 = {{1{spriteYPositionReg_0[9]}},spriteYPositionReg_0}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_432 = $signed(_T_431) - $signed(_GEN_1120); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_436 = $signed(inSpriteX_0) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_437 = $signed(inSpriteX_0) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_438 = _T_436 & _T_437; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_0 = _T_432[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_439 = $signed(inSpriteY_0) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_440 = _T_438 & _T_439; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_441 = $signed(inSpriteY_0) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_1 = $signed(_T_425) - $signed(spriteXPositionReg_1); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1122 = {{1{spriteYPositionReg_1[9]}},spriteYPositionReg_1}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_451 = $signed(_T_431) - $signed(_GEN_1122); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_455 = $signed(inSpriteX_1) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_456 = $signed(inSpriteX_1) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_457 = _T_455 & _T_456; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_1 = _T_451[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_458 = $signed(inSpriteY_1) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_459 = _T_457 & _T_458; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_460 = $signed(inSpriteY_1) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_2 = $signed(_T_425) - $signed(spriteXPositionReg_2); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1124 = {{1{spriteYPositionReg_2[9]}},spriteYPositionReg_2}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_470 = $signed(_T_431) - $signed(_GEN_1124); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_474 = $signed(inSpriteX_2) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_475 = $signed(inSpriteX_2) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_476 = _T_474 & _T_475; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_2 = _T_470[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_477 = $signed(inSpriteY_2) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_478 = _T_476 & _T_477; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_479 = $signed(inSpriteY_2) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_3 = $signed(_T_425) - $signed(spriteXPositionReg_3); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1126 = {{1{spriteYPositionReg_3[9]}},spriteYPositionReg_3}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_489 = $signed(_T_431) - $signed(_GEN_1126); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_493 = $signed(inSpriteX_3) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_494 = $signed(inSpriteX_3) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_495 = _T_493 & _T_494; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_3 = _T_489[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_496 = $signed(inSpriteY_3) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_497 = _T_495 & _T_496; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_498 = $signed(inSpriteY_3) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_4 = $signed(_T_425) - $signed(spriteXPositionReg_4); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1128 = {{1{spriteYPositionReg_4[9]}},spriteYPositionReg_4}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_508 = $signed(_T_431) - $signed(_GEN_1128); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_512 = $signed(inSpriteX_4) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_513 = $signed(inSpriteX_4) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_514 = _T_512 & _T_513; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_4 = _T_508[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_515 = $signed(inSpriteY_4) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_516 = _T_514 & _T_515; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_517 = $signed(inSpriteY_4) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_5 = $signed(_T_425) - $signed(spriteXPositionReg_5); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1130 = {{1{spriteYPositionReg_5[9]}},spriteYPositionReg_5}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_527 = $signed(_T_431) - $signed(_GEN_1130); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_531 = $signed(inSpriteX_5) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_532 = $signed(inSpriteX_5) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_533 = _T_531 & _T_532; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_5 = _T_527[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_534 = $signed(inSpriteY_5) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_535 = _T_533 & _T_534; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_536 = $signed(inSpriteY_5) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_6 = $signed(_T_425) - $signed(spriteXPositionReg_6); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1132 = {{1{spriteYPositionReg_6[9]}},spriteYPositionReg_6}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_546 = $signed(_T_431) - $signed(_GEN_1132); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_550 = $signed(inSpriteX_6) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_551 = $signed(inSpriteX_6) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_552 = _T_550 & _T_551; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_6 = _T_546[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_553 = $signed(inSpriteY_6) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_554 = _T_552 & _T_553; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_555 = $signed(inSpriteY_6) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_7 = $signed(_T_425) - $signed(spriteXPositionReg_7); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1134 = {{1{spriteYPositionReg_7[9]}},spriteYPositionReg_7}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_565 = $signed(_T_431) - $signed(_GEN_1134); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_569 = $signed(inSpriteX_7) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_570 = $signed(inSpriteX_7) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_571 = _T_569 & _T_570; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_7 = _T_565[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_572 = $signed(inSpriteY_7) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_573 = _T_571 & _T_572; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_574 = $signed(inSpriteY_7) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_8 = $signed(_T_425) - $signed(spriteXPositionReg_8); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1136 = {{1{spriteYPositionReg_8[9]}},spriteYPositionReg_8}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_584 = $signed(_T_431) - $signed(_GEN_1136); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_588 = $signed(inSpriteX_8) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_589 = $signed(inSpriteX_8) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_590 = _T_588 & _T_589; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_8 = _T_584[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_591 = $signed(inSpriteY_8) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_592 = _T_590 & _T_591; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_593 = $signed(inSpriteY_8) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_9 = $signed(_T_425) - $signed(spriteXPositionReg_9); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1138 = {{1{spriteYPositionReg_9[9]}},spriteYPositionReg_9}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_603 = $signed(_T_431) - $signed(_GEN_1138); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_607 = $signed(inSpriteX_9) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_608 = $signed(inSpriteX_9) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_609 = _T_607 & _T_608; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_9 = _T_603[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_610 = $signed(inSpriteY_9) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_611 = _T_609 & _T_610; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_612 = $signed(inSpriteY_9) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_10 = $signed(_T_425) - $signed(spriteXPositionReg_10); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1140 = {{1{spriteYPositionReg_10[9]}},spriteYPositionReg_10}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_622 = $signed(_T_431) - $signed(_GEN_1140); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_626 = $signed(inSpriteX_10) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_627 = $signed(inSpriteX_10) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_628 = _T_626 & _T_627; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_10 = _T_622[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_629 = $signed(inSpriteY_10) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_630 = _T_628 & _T_629; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_631 = $signed(inSpriteY_10) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_11 = $signed(_T_425) - $signed(spriteXPositionReg_11); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1142 = {{1{spriteYPositionReg_11[9]}},spriteYPositionReg_11}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_641 = $signed(_T_431) - $signed(_GEN_1142); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_645 = $signed(inSpriteX_11) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_646 = $signed(inSpriteX_11) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_647 = _T_645 & _T_646; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_11 = _T_641[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_648 = $signed(inSpriteY_11) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_649 = _T_647 & _T_648; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_650 = $signed(inSpriteY_11) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_12 = $signed(_T_425) - $signed(spriteXPositionReg_12); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1144 = {{1{spriteYPositionReg_12[9]}},spriteYPositionReg_12}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_660 = $signed(_T_431) - $signed(_GEN_1144); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_664 = $signed(inSpriteX_12) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_665 = $signed(inSpriteX_12) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_666 = _T_664 & _T_665; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_12 = _T_660[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_667 = $signed(inSpriteY_12) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_668 = _T_666 & _T_667; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_669 = $signed(inSpriteY_12) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_13 = $signed(_T_425) - $signed(spriteXPositionReg_13); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1146 = {{1{spriteYPositionReg_13[9]}},spriteYPositionReg_13}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_679 = $signed(_T_431) - $signed(_GEN_1146); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_683 = $signed(inSpriteX_13) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_684 = $signed(inSpriteX_13) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_685 = _T_683 & _T_684; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_13 = _T_679[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_686 = $signed(inSpriteY_13) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_687 = _T_685 & _T_686; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_688 = $signed(inSpriteY_13) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_14 = $signed(_T_425) - $signed(spriteXPositionReg_14); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1148 = {{1{spriteYPositionReg_14[9]}},spriteYPositionReg_14}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_698 = $signed(_T_431) - $signed(_GEN_1148); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_702 = $signed(inSpriteX_14) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_703 = $signed(inSpriteX_14) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_704 = _T_702 & _T_703; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_14 = _T_698[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_705 = $signed(inSpriteY_14) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_706 = _T_704 & _T_705; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_707 = $signed(inSpriteY_14) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_15 = $signed(_T_425) - $signed(spriteXPositionReg_15); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1150 = {{1{spriteYPositionReg_15[9]}},spriteYPositionReg_15}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_717 = $signed(_T_431) - $signed(_GEN_1150); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_721 = $signed(inSpriteX_15) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_722 = $signed(inSpriteX_15) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_723 = _T_721 & _T_722; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_15 = _T_717[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_724 = $signed(inSpriteY_15) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_725 = _T_723 & _T_724; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_726 = $signed(inSpriteY_15) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_16 = $signed(_T_425) - $signed(spriteXPositionReg_16); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1152 = {{1{spriteYPositionReg_16[9]}},spriteYPositionReg_16}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_736 = $signed(_T_431) - $signed(_GEN_1152); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_740 = $signed(inSpriteX_16) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_741 = $signed(inSpriteX_16) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_742 = _T_740 & _T_741; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_16 = _T_736[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_743 = $signed(inSpriteY_16) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_744 = _T_742 & _T_743; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_745 = $signed(inSpriteY_16) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_17 = $signed(_T_425) - $signed(spriteXPositionReg_17); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1154 = {{1{spriteYPositionReg_17[9]}},spriteYPositionReg_17}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_755 = $signed(_T_431) - $signed(_GEN_1154); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_759 = $signed(inSpriteX_17) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_760 = $signed(inSpriteX_17) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_761 = _T_759 & _T_760; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_17 = _T_755[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_762 = $signed(inSpriteY_17) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_763 = _T_761 & _T_762; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_764 = $signed(inSpriteY_17) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_18 = $signed(_T_425) - $signed(spriteXPositionReg_18); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1156 = {{1{spriteYPositionReg_18[9]}},spriteYPositionReg_18}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_774 = $signed(_T_431) - $signed(_GEN_1156); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_778 = $signed(inSpriteX_18) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_779 = $signed(inSpriteX_18) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_780 = _T_778 & _T_779; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_18 = _T_774[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_781 = $signed(inSpriteY_18) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_782 = _T_780 & _T_781; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_783 = $signed(inSpriteY_18) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_19 = $signed(_T_425) - $signed(spriteXPositionReg_19); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1158 = {{1{spriteYPositionReg_19[9]}},spriteYPositionReg_19}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_793 = $signed(_T_431) - $signed(_GEN_1158); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_797 = $signed(inSpriteX_19) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_798 = $signed(inSpriteX_19) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_799 = _T_797 & _T_798; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_19 = _T_793[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_800 = $signed(inSpriteY_19) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_801 = _T_799 & _T_800; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_802 = $signed(inSpriteY_19) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_20 = $signed(_T_425) - $signed(spriteXPositionReg_20); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1160 = {{1{spriteYPositionReg_20[9]}},spriteYPositionReg_20}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_812 = $signed(_T_431) - $signed(_GEN_1160); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_816 = $signed(inSpriteX_20) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_817 = $signed(inSpriteX_20) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_818 = _T_816 & _T_817; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_20 = _T_812[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_819 = $signed(inSpriteY_20) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_820 = _T_818 & _T_819; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_821 = $signed(inSpriteY_20) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_21 = $signed(_T_425) - $signed(spriteXPositionReg_21); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1162 = {{1{spriteYPositionReg_21[9]}},spriteYPositionReg_21}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_831 = $signed(_T_431) - $signed(_GEN_1162); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_835 = $signed(inSpriteX_21) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_836 = $signed(inSpriteX_21) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_837 = _T_835 & _T_836; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_21 = _T_831[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_838 = $signed(inSpriteY_21) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_839 = _T_837 & _T_838; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_840 = $signed(inSpriteY_21) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_22 = $signed(_T_425) - $signed(spriteXPositionReg_22); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1164 = {{1{spriteYPositionReg_22[9]}},spriteYPositionReg_22}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_850 = $signed(_T_431) - $signed(_GEN_1164); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_854 = $signed(inSpriteX_22) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_855 = $signed(inSpriteX_22) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_856 = _T_854 & _T_855; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_22 = _T_850[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_857 = $signed(inSpriteY_22) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_858 = _T_856 & _T_857; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_859 = $signed(inSpriteY_22) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_23 = $signed(_T_425) - $signed(spriteXPositionReg_23); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1166 = {{1{spriteYPositionReg_23[9]}},spriteYPositionReg_23}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_869 = $signed(_T_431) - $signed(_GEN_1166); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_873 = $signed(inSpriteX_23) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_874 = $signed(inSpriteX_23) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_875 = _T_873 & _T_874; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_23 = _T_869[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_876 = $signed(inSpriteY_23) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_877 = _T_875 & _T_876; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_878 = $signed(inSpriteY_23) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_24 = $signed(_T_425) - $signed(spriteXPositionReg_24); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1168 = {{1{spriteYPositionReg_24[9]}},spriteYPositionReg_24}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_888 = $signed(_T_431) - $signed(_GEN_1168); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_892 = $signed(inSpriteX_24) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_893 = $signed(inSpriteX_24) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_894 = _T_892 & _T_893; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_24 = _T_888[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_895 = $signed(inSpriteY_24) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_896 = _T_894 & _T_895; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_897 = $signed(inSpriteY_24) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_25 = $signed(_T_425) - $signed(spriteXPositionReg_25); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1170 = {{1{spriteYPositionReg_25[9]}},spriteYPositionReg_25}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_907 = $signed(_T_431) - $signed(_GEN_1170); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_911 = $signed(inSpriteX_25) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_912 = $signed(inSpriteX_25) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_913 = _T_911 & _T_912; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_25 = _T_907[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_914 = $signed(inSpriteY_25) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_915 = _T_913 & _T_914; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_916 = $signed(inSpriteY_25) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_26 = $signed(_T_425) - $signed(spriteXPositionReg_26); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1172 = {{1{spriteYPositionReg_26[9]}},spriteYPositionReg_26}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_926 = $signed(_T_431) - $signed(_GEN_1172); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_930 = $signed(inSpriteX_26) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_931 = $signed(inSpriteX_26) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_932 = _T_930 & _T_931; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_26 = _T_926[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_933 = $signed(inSpriteY_26) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_934 = _T_932 & _T_933; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_935 = $signed(inSpriteY_26) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_27 = $signed(_T_425) - $signed(spriteXPositionReg_27); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1174 = {{1{spriteYPositionReg_27[9]}},spriteYPositionReg_27}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_945 = $signed(_T_431) - $signed(_GEN_1174); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_949 = $signed(inSpriteX_27) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_950 = $signed(inSpriteX_27) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_951 = _T_949 & _T_950; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_27 = _T_945[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_952 = $signed(inSpriteY_27) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_953 = _T_951 & _T_952; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_954 = $signed(inSpriteY_27) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_28 = $signed(_T_425) - $signed(spriteXPositionReg_28); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1176 = {{1{spriteYPositionReg_28[9]}},spriteYPositionReg_28}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_964 = $signed(_T_431) - $signed(_GEN_1176); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_968 = $signed(inSpriteX_28) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_969 = $signed(inSpriteX_28) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_970 = _T_968 & _T_969; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_28 = _T_964[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_971 = $signed(inSpriteY_28) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_972 = _T_970 & _T_971; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_973 = $signed(inSpriteY_28) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_29 = $signed(_T_425) - $signed(spriteXPositionReg_29); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1178 = {{1{spriteYPositionReg_29[9]}},spriteYPositionReg_29}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_983 = $signed(_T_431) - $signed(_GEN_1178); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_987 = $signed(inSpriteX_29) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_988 = $signed(inSpriteX_29) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_989 = _T_987 & _T_988; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_29 = _T_983[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_990 = $signed(inSpriteY_29) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_991 = _T_989 & _T_990; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_992 = $signed(inSpriteY_29) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_30 = $signed(_T_425) - $signed(spriteXPositionReg_30); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1180 = {{1{spriteYPositionReg_30[9]}},spriteYPositionReg_30}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1002 = $signed(_T_431) - $signed(_GEN_1180); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1006 = $signed(inSpriteX_30) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1007 = $signed(inSpriteX_30) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1008 = _T_1006 & _T_1007; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_30 = _T_1002[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1009 = $signed(inSpriteY_30) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1010 = _T_1008 & _T_1009; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1011 = $signed(inSpriteY_30) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_31 = $signed(_T_425) - $signed(spriteXPositionReg_31); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1182 = {{1{spriteYPositionReg_31[9]}},spriteYPositionReg_31}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1021 = $signed(_T_431) - $signed(_GEN_1182); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1025 = $signed(inSpriteX_31) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1026 = $signed(inSpriteX_31) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1027 = _T_1025 & _T_1026; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_31 = _T_1021[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1028 = $signed(inSpriteY_31) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1029 = _T_1027 & _T_1028; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1030 = $signed(inSpriteY_31) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_32 = $signed(_T_425) - $signed(spriteXPositionReg_32); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1184 = {{1{spriteYPositionReg_32[9]}},spriteYPositionReg_32}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1040 = $signed(_T_431) - $signed(_GEN_1184); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1044 = $signed(inSpriteX_32) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1045 = $signed(inSpriteX_32) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1046 = _T_1044 & _T_1045; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_32 = _T_1040[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1047 = $signed(inSpriteY_32) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1048 = _T_1046 & _T_1047; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1049 = $signed(inSpriteY_32) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_33 = $signed(_T_425) - $signed(spriteXPositionReg_33); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1186 = {{1{spriteYPositionReg_33[9]}},spriteYPositionReg_33}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1059 = $signed(_T_431) - $signed(_GEN_1186); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1063 = $signed(inSpriteX_33) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1064 = $signed(inSpriteX_33) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1065 = _T_1063 & _T_1064; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_33 = _T_1059[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1066 = $signed(inSpriteY_33) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1067 = _T_1065 & _T_1066; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1068 = $signed(inSpriteY_33) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_34 = $signed(_T_425) - $signed(spriteXPositionReg_34); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1188 = {{1{spriteYPositionReg_34[9]}},spriteYPositionReg_34}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1078 = $signed(_T_431) - $signed(_GEN_1188); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1082 = $signed(inSpriteX_34) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1083 = $signed(inSpriteX_34) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1084 = _T_1082 & _T_1083; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_34 = _T_1078[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1085 = $signed(inSpriteY_34) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1086 = _T_1084 & _T_1085; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1087 = $signed(inSpriteY_34) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_35 = $signed(_T_425) - $signed(spriteXPositionReg_35); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1190 = {{1{spriteYPositionReg_35[9]}},spriteYPositionReg_35}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1097 = $signed(_T_431) - $signed(_GEN_1190); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1101 = $signed(inSpriteX_35) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1102 = $signed(inSpriteX_35) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1103 = _T_1101 & _T_1102; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_35 = _T_1097[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1104 = $signed(inSpriteY_35) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1105 = _T_1103 & _T_1104; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1106 = $signed(inSpriteY_35) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_36 = $signed(_T_425) - $signed(spriteXPositionReg_36); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1192 = {{1{spriteYPositionReg_36[9]}},spriteYPositionReg_36}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1116 = $signed(_T_431) - $signed(_GEN_1192); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1120 = $signed(inSpriteX_36) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1121 = $signed(inSpriteX_36) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1122 = _T_1120 & _T_1121; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_36 = _T_1116[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1123 = $signed(inSpriteY_36) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1124 = _T_1122 & _T_1123; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1125 = $signed(inSpriteY_36) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_37 = $signed(_T_425) - $signed(spriteXPositionReg_37); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1194 = {{1{spriteYPositionReg_37[9]}},spriteYPositionReg_37}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1135 = $signed(_T_431) - $signed(_GEN_1194); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1139 = $signed(inSpriteX_37) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1140 = $signed(inSpriteX_37) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1141 = _T_1139 & _T_1140; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_37 = _T_1135[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1142 = $signed(inSpriteY_37) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1143 = _T_1141 & _T_1142; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1144 = $signed(inSpriteY_37) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_38 = $signed(_T_425) - $signed(spriteXPositionReg_38); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1196 = {{1{spriteYPositionReg_38[9]}},spriteYPositionReg_38}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1154 = $signed(_T_431) - $signed(_GEN_1196); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1158 = $signed(inSpriteX_38) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1159 = $signed(inSpriteX_38) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1160 = _T_1158 & _T_1159; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_38 = _T_1154[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1161 = $signed(inSpriteY_38) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1162 = _T_1160 & _T_1161; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1163 = $signed(inSpriteY_38) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_39 = $signed(_T_425) - $signed(spriteXPositionReg_39); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1198 = {{1{spriteYPositionReg_39[9]}},spriteYPositionReg_39}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1173 = $signed(_T_431) - $signed(_GEN_1198); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1177 = $signed(inSpriteX_39) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1178 = $signed(inSpriteX_39) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1179 = _T_1177 & _T_1178; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_39 = _T_1173[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1180 = $signed(inSpriteY_39) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1181 = _T_1179 & _T_1180; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1182 = $signed(inSpriteY_39) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_40 = $signed(_T_425) - $signed(spriteXPositionReg_40); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1200 = {{1{spriteYPositionReg_40[9]}},spriteYPositionReg_40}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1192 = $signed(_T_431) - $signed(_GEN_1200); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1196 = $signed(inSpriteX_40) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1197 = $signed(inSpriteX_40) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1198 = _T_1196 & _T_1197; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_40 = _T_1192[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1199 = $signed(inSpriteY_40) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1200 = _T_1198 & _T_1199; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1201 = $signed(inSpriteY_40) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_41 = $signed(_T_425) - $signed(spriteXPositionReg_41); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1202 = {{1{spriteYPositionReg_41[9]}},spriteYPositionReg_41}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1211 = $signed(_T_431) - $signed(_GEN_1202); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1215 = $signed(inSpriteX_41) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1216 = $signed(inSpriteX_41) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1217 = _T_1215 & _T_1216; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_41 = _T_1211[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1218 = $signed(inSpriteY_41) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1219 = _T_1217 & _T_1218; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1220 = $signed(inSpriteY_41) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_42 = $signed(_T_425) - $signed(spriteXPositionReg_42); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1204 = {{1{spriteYPositionReg_42[9]}},spriteYPositionReg_42}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1230 = $signed(_T_431) - $signed(_GEN_1204); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1234 = $signed(inSpriteX_42) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1235 = $signed(inSpriteX_42) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1236 = _T_1234 & _T_1235; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_42 = _T_1230[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1237 = $signed(inSpriteY_42) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1238 = _T_1236 & _T_1237; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1239 = $signed(inSpriteY_42) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_43 = $signed(_T_425) - $signed(spriteXPositionReg_43); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1206 = {{1{spriteYPositionReg_43[9]}},spriteYPositionReg_43}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1249 = $signed(_T_431) - $signed(_GEN_1206); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1253 = $signed(inSpriteX_43) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1254 = $signed(inSpriteX_43) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1255 = _T_1253 & _T_1254; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_43 = _T_1249[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1256 = $signed(inSpriteY_43) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1257 = _T_1255 & _T_1256; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1258 = $signed(inSpriteY_43) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_44 = $signed(_T_425) - $signed(spriteXPositionReg_44); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1208 = {{1{spriteYPositionReg_44[9]}},spriteYPositionReg_44}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1268 = $signed(_T_431) - $signed(_GEN_1208); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1272 = $signed(inSpriteX_44) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1273 = $signed(inSpriteX_44) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1274 = _T_1272 & _T_1273; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_44 = _T_1268[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1275 = $signed(inSpriteY_44) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1276 = _T_1274 & _T_1275; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1277 = $signed(inSpriteY_44) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_45 = $signed(_T_425) - $signed(spriteXPositionReg_45); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1210 = {{1{spriteYPositionReg_45[9]}},spriteYPositionReg_45}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1287 = $signed(_T_431) - $signed(_GEN_1210); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1291 = $signed(inSpriteX_45) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1292 = $signed(inSpriteX_45) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1293 = _T_1291 & _T_1292; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_45 = _T_1287[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1294 = $signed(inSpriteY_45) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1295 = _T_1293 & _T_1294; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1296 = $signed(inSpriteY_45) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_46 = $signed(_T_425) - $signed(spriteXPositionReg_46); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1212 = {{1{spriteYPositionReg_46[9]}},spriteYPositionReg_46}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1306 = $signed(_T_431) - $signed(_GEN_1212); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1310 = $signed(inSpriteX_46) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1311 = $signed(inSpriteX_46) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1312 = _T_1310 & _T_1311; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_46 = _T_1306[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1313 = $signed(inSpriteY_46) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1314 = _T_1312 & _T_1313; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1315 = $signed(inSpriteY_46) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_47 = $signed(_T_425) - $signed(spriteXPositionReg_47); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1214 = {{1{spriteYPositionReg_47[9]}},spriteYPositionReg_47}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1325 = $signed(_T_431) - $signed(_GEN_1214); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1329 = $signed(inSpriteX_47) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1330 = $signed(inSpriteX_47) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1331 = _T_1329 & _T_1330; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_47 = _T_1325[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1332 = $signed(inSpriteY_47) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1333 = _T_1331 & _T_1332; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1334 = $signed(inSpriteY_47) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_48 = $signed(_T_425) - $signed(spriteXPositionReg_48); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1216 = {{1{spriteYPositionReg_48[9]}},spriteYPositionReg_48}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1344 = $signed(_T_431) - $signed(_GEN_1216); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1348 = $signed(inSpriteX_48) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1349 = $signed(inSpriteX_48) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1350 = _T_1348 & _T_1349; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_48 = _T_1344[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1351 = $signed(inSpriteY_48) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1352 = _T_1350 & _T_1351; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1353 = $signed(inSpriteY_48) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_49 = $signed(_T_425) - $signed(spriteXPositionReg_49); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1218 = {{1{spriteYPositionReg_49[9]}},spriteYPositionReg_49}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1363 = $signed(_T_431) - $signed(_GEN_1218); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1367 = $signed(inSpriteX_49) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1368 = $signed(inSpriteX_49) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1369 = _T_1367 & _T_1368; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_49 = _T_1363[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1370 = $signed(inSpriteY_49) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1371 = _T_1369 & _T_1370; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1372 = $signed(inSpriteY_49) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_50 = $signed(_T_425) - $signed(spriteXPositionReg_50); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1220 = {{1{spriteYPositionReg_50[9]}},spriteYPositionReg_50}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1382 = $signed(_T_431) - $signed(_GEN_1220); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1386 = $signed(inSpriteX_50) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1387 = $signed(inSpriteX_50) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1388 = _T_1386 & _T_1387; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_50 = _T_1382[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1389 = $signed(inSpriteY_50) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1390 = _T_1388 & _T_1389; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1391 = $signed(inSpriteY_50) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_51 = $signed(_T_425) - $signed(spriteXPositionReg_51); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1222 = {{1{spriteYPositionReg_51[9]}},spriteYPositionReg_51}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1401 = $signed(_T_431) - $signed(_GEN_1222); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1405 = $signed(inSpriteX_51) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1406 = $signed(inSpriteX_51) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1407 = _T_1405 & _T_1406; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_51 = _T_1401[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1408 = $signed(inSpriteY_51) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1409 = _T_1407 & _T_1408; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1410 = $signed(inSpriteY_51) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_52 = $signed(_T_425) - $signed(spriteXPositionReg_52); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1224 = {{1{spriteYPositionReg_52[9]}},spriteYPositionReg_52}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1420 = $signed(_T_431) - $signed(_GEN_1224); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1424 = $signed(inSpriteX_52) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1425 = $signed(inSpriteX_52) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1426 = _T_1424 & _T_1425; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_52 = _T_1420[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1427 = $signed(inSpriteY_52) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1428 = _T_1426 & _T_1427; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1429 = $signed(inSpriteY_52) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_53 = $signed(_T_425) - $signed(spriteXPositionReg_53); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1226 = {{1{spriteYPositionReg_53[9]}},spriteYPositionReg_53}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1439 = $signed(_T_431) - $signed(_GEN_1226); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1443 = $signed(inSpriteX_53) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1444 = $signed(inSpriteX_53) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1445 = _T_1443 & _T_1444; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_53 = _T_1439[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1446 = $signed(inSpriteY_53) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1447 = _T_1445 & _T_1446; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1448 = $signed(inSpriteY_53) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_54 = $signed(_T_425) - $signed(spriteXPositionReg_54); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1228 = {{1{spriteYPositionReg_54[9]}},spriteYPositionReg_54}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1458 = $signed(_T_431) - $signed(_GEN_1228); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1462 = $signed(inSpriteX_54) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1463 = $signed(inSpriteX_54) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1464 = _T_1462 & _T_1463; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_54 = _T_1458[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1465 = $signed(inSpriteY_54) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1466 = _T_1464 & _T_1465; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1467 = $signed(inSpriteY_54) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_55 = $signed(_T_425) - $signed(spriteXPositionReg_55); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1230 = {{1{spriteYPositionReg_55[9]}},spriteYPositionReg_55}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1477 = $signed(_T_431) - $signed(_GEN_1230); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1481 = $signed(inSpriteX_55) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1482 = $signed(inSpriteX_55) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1483 = _T_1481 & _T_1482; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_55 = _T_1477[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1484 = $signed(inSpriteY_55) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1485 = _T_1483 & _T_1484; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1486 = $signed(inSpriteY_55) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_56 = $signed(_T_425) - $signed(spriteXPositionReg_56); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1232 = {{1{spriteYPositionReg_56[9]}},spriteYPositionReg_56}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1496 = $signed(_T_431) - $signed(_GEN_1232); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1500 = $signed(inSpriteX_56) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1501 = $signed(inSpriteX_56) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1502 = _T_1500 & _T_1501; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_56 = _T_1496[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1503 = $signed(inSpriteY_56) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1504 = _T_1502 & _T_1503; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1505 = $signed(inSpriteY_56) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_57 = $signed(_T_425) - $signed(spriteXPositionReg_57); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1234 = {{1{spriteYPositionReg_57[9]}},spriteYPositionReg_57}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1515 = $signed(_T_431) - $signed(_GEN_1234); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1519 = $signed(inSpriteX_57) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1520 = $signed(inSpriteX_57) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1521 = _T_1519 & _T_1520; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_57 = _T_1515[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1522 = $signed(inSpriteY_57) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1523 = _T_1521 & _T_1522; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1524 = $signed(inSpriteY_57) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_58 = $signed(_T_425) - $signed(spriteXPositionReg_58); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1236 = {{1{spriteYPositionReg_58[9]}},spriteYPositionReg_58}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1534 = $signed(_T_431) - $signed(_GEN_1236); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1538 = $signed(inSpriteX_58) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1539 = $signed(inSpriteX_58) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1540 = _T_1538 & _T_1539; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_58 = _T_1534[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1541 = $signed(inSpriteY_58) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1542 = _T_1540 & _T_1541; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1543 = $signed(inSpriteY_58) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_59 = $signed(_T_425) - $signed(spriteXPositionReg_59); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1238 = {{1{spriteYPositionReg_59[9]}},spriteYPositionReg_59}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1553 = $signed(_T_431) - $signed(_GEN_1238); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1557 = $signed(inSpriteX_59) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1558 = $signed(inSpriteX_59) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1559 = _T_1557 & _T_1558; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_59 = _T_1553[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1560 = $signed(inSpriteY_59) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1561 = _T_1559 & _T_1560; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1562 = $signed(inSpriteY_59) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_60 = $signed(_T_425) - $signed(spriteXPositionReg_60); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1240 = {{1{spriteYPositionReg_60[9]}},spriteYPositionReg_60}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1572 = $signed(_T_431) - $signed(_GEN_1240); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1576 = $signed(inSpriteX_60) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1577 = $signed(inSpriteX_60) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1578 = _T_1576 & _T_1577; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_60 = _T_1572[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1579 = $signed(inSpriteY_60) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1580 = _T_1578 & _T_1579; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1581 = $signed(inSpriteY_60) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_61 = $signed(_T_425) - $signed(spriteXPositionReg_61); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1242 = {{1{spriteYPositionReg_61[9]}},spriteYPositionReg_61}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1591 = $signed(_T_431) - $signed(_GEN_1242); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1595 = $signed(inSpriteX_61) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1596 = $signed(inSpriteX_61) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1597 = _T_1595 & _T_1596; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_61 = _T_1591[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1598 = $signed(inSpriteY_61) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1599 = _T_1597 & _T_1598; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1600 = $signed(inSpriteY_61) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_62 = $signed(_T_425) - $signed(spriteXPositionReg_62); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1244 = {{1{spriteYPositionReg_62[9]}},spriteYPositionReg_62}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1610 = $signed(_T_431) - $signed(_GEN_1244); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1614 = $signed(inSpriteX_62) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1615 = $signed(inSpriteX_62) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1616 = _T_1614 & _T_1615; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_62 = _T_1610[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1617 = $signed(inSpriteY_62) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1618 = _T_1616 & _T_1617; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1619 = $signed(inSpriteY_62) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_63 = $signed(_T_425) - $signed(spriteXPositionReg_63); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1246 = {{1{spriteYPositionReg_63[9]}},spriteYPositionReg_63}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1629 = $signed(_T_431) - $signed(_GEN_1246); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1633 = $signed(inSpriteX_63) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1634 = $signed(inSpriteX_63) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1635 = _T_1633 & _T_1634; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_63 = _T_1629[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1636 = $signed(inSpriteY_63) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1637 = _T_1635 & _T_1636; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1638 = $signed(inSpriteY_63) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_64 = $signed(_T_425) - $signed(spriteXPositionReg_64); // @[GraphicEngineVGA.scala 281:54]
  wire [11:0] _T_1648 = $signed(_T_431) - 11'sh0; // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1652 = $signed(inSpriteX_64) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1653 = $signed(inSpriteX_64) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1654 = _T_1652 & _T_1653; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_64 = _T_1648[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1655 = $signed(inSpriteY_64) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1656 = _T_1654 & _T_1655; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1657 = $signed(inSpriteY_64) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_65 = $signed(_T_425) - $signed(spriteXPositionReg_65); // @[GraphicEngineVGA.scala 281:54]
  wire  _T_1671 = $signed(inSpriteX_65) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1672 = $signed(inSpriteX_65) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1673 = _T_1671 & _T_1672; // @[GraphicEngineVGA.scala 293:40]
  wire  _T_1675 = _T_1673 & _T_1655; // @[GraphicEngineVGA.scala 293:63]
  wire [11:0] inSpriteX_66 = $signed(_T_425) - $signed(spriteXPositionReg_66); // @[GraphicEngineVGA.scala 281:54]
  wire  _T_1690 = $signed(inSpriteX_66) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1691 = $signed(inSpriteX_66) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1692 = _T_1690 & _T_1691; // @[GraphicEngineVGA.scala 293:40]
  wire  _T_1694 = _T_1692 & _T_1655; // @[GraphicEngineVGA.scala 293:63]
  wire [11:0] inSpriteX_67 = $signed(_T_425) - $signed(spriteXPositionReg_67); // @[GraphicEngineVGA.scala 281:54]
  wire  _T_1709 = $signed(inSpriteX_67) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1710 = $signed(inSpriteX_67) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1711 = _T_1709 & _T_1710; // @[GraphicEngineVGA.scala 293:40]
  wire  _T_1713 = _T_1711 & _T_1655; // @[GraphicEngineVGA.scala 293:63]
  wire [11:0] inSpriteX_68 = $signed(_T_425) - $signed(spriteXPositionReg_68); // @[GraphicEngineVGA.scala 281:54]
  wire  _T_1728 = $signed(inSpriteX_68) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1729 = $signed(inSpriteX_68) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1730 = _T_1728 & _T_1729; // @[GraphicEngineVGA.scala 293:40]
  wire  _T_1732 = _T_1730 & _T_1655; // @[GraphicEngineVGA.scala 293:63]
  wire [11:0] inSpriteX_69 = $signed(_T_425) - $signed(spriteXPositionReg_69); // @[GraphicEngineVGA.scala 281:54]
  wire  _T_1747 = $signed(inSpriteX_69) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1748 = $signed(inSpriteX_69) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1749 = _T_1747 & _T_1748; // @[GraphicEngineVGA.scala 293:40]
  wire  _T_1751 = _T_1749 & _T_1655; // @[GraphicEngineVGA.scala 293:63]
  wire [11:0] inSpriteX_70 = $signed(_T_425) - $signed(spriteXPositionReg_70); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1254 = {{1{spriteYPositionReg_70[9]}},spriteYPositionReg_70}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1762 = $signed(_T_431) - $signed(_GEN_1254); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1766 = $signed(inSpriteX_70) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1767 = $signed(inSpriteX_70) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1768 = _T_1766 & _T_1767; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_70 = _T_1762[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1769 = $signed(inSpriteY_70) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1770 = _T_1768 & _T_1769; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1771 = $signed(inSpriteY_70) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_71 = $signed(_T_425) - $signed(spriteXPositionReg_71); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1256 = {{1{spriteYPositionReg_71[9]}},spriteYPositionReg_71}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1781 = $signed(_T_431) - $signed(_GEN_1256); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1785 = $signed(inSpriteX_71) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1786 = $signed(inSpriteX_71) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1787 = _T_1785 & _T_1786; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_71 = _T_1781[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1788 = $signed(inSpriteY_71) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1789 = _T_1787 & _T_1788; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1790 = $signed(inSpriteY_71) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_72 = $signed(_T_425) - $signed(spriteXPositionReg_72); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1258 = {{1{spriteYPositionReg_72[9]}},spriteYPositionReg_72}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1800 = $signed(_T_431) - $signed(_GEN_1258); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1804 = $signed(inSpriteX_72) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1805 = $signed(inSpriteX_72) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1806 = _T_1804 & _T_1805; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_72 = _T_1800[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1807 = $signed(inSpriteY_72) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1808 = _T_1806 & _T_1807; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1809 = $signed(inSpriteY_72) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_73 = $signed(_T_425) - $signed(spriteXPositionReg_73); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1260 = {{1{spriteYPositionReg_73[9]}},spriteYPositionReg_73}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1819 = $signed(_T_431) - $signed(_GEN_1260); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1823 = $signed(inSpriteX_73) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1824 = $signed(inSpriteX_73) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1825 = _T_1823 & _T_1824; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_73 = _T_1819[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1826 = $signed(inSpriteY_73) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1827 = _T_1825 & _T_1826; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1828 = $signed(inSpriteY_73) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_74 = $signed(_T_425) - $signed(spriteXPositionReg_74); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1262 = {{1{spriteYPositionReg_74[9]}},spriteYPositionReg_74}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1838 = $signed(_T_431) - $signed(_GEN_1262); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1842 = $signed(inSpriteX_74) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1843 = $signed(inSpriteX_74) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1844 = _T_1842 & _T_1843; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_74 = _T_1838[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1845 = $signed(inSpriteY_74) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1846 = _T_1844 & _T_1845; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1847 = $signed(inSpriteY_74) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_75 = $signed(_T_425) - $signed(spriteXPositionReg_75); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1264 = {{1{spriteYPositionReg_75[9]}},spriteYPositionReg_75}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1857 = $signed(_T_431) - $signed(_GEN_1264); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1861 = $signed(inSpriteX_75) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1862 = $signed(inSpriteX_75) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1863 = _T_1861 & _T_1862; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_75 = _T_1857[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1864 = $signed(inSpriteY_75) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1865 = _T_1863 & _T_1864; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1866 = $signed(inSpriteY_75) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_76 = $signed(_T_425) - $signed(spriteXPositionReg_76); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1266 = {{1{spriteYPositionReg_76[9]}},spriteYPositionReg_76}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1876 = $signed(_T_431) - $signed(_GEN_1266); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1880 = $signed(inSpriteX_76) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1881 = $signed(inSpriteX_76) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1882 = _T_1880 & _T_1881; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_76 = _T_1876[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1883 = $signed(inSpriteY_76) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1884 = _T_1882 & _T_1883; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1885 = $signed(inSpriteY_76) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_77 = $signed(_T_425) - $signed(spriteXPositionReg_77); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1268 = {{1{spriteYPositionReg_77[9]}},spriteYPositionReg_77}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1895 = $signed(_T_431) - $signed(_GEN_1268); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1899 = $signed(inSpriteX_77) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1900 = $signed(inSpriteX_77) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1901 = _T_1899 & _T_1900; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_77 = _T_1895[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1902 = $signed(inSpriteY_77) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1903 = _T_1901 & _T_1902; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1904 = $signed(inSpriteY_77) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_78 = $signed(_T_425) - $signed(spriteXPositionReg_78); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1270 = {{1{spriteYPositionReg_78[9]}},spriteYPositionReg_78}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1914 = $signed(_T_431) - $signed(_GEN_1270); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1918 = $signed(inSpriteX_78) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1919 = $signed(inSpriteX_78) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1920 = _T_1918 & _T_1919; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_78 = _T_1914[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1921 = $signed(inSpriteY_78) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1922 = _T_1920 & _T_1921; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1923 = $signed(inSpriteY_78) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_79 = $signed(_T_425) - $signed(spriteXPositionReg_79); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1272 = {{1{spriteYPositionReg_79[9]}},spriteYPositionReg_79}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1933 = $signed(_T_431) - $signed(_GEN_1272); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1937 = $signed(inSpriteX_79) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1938 = $signed(inSpriteX_79) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1939 = _T_1937 & _T_1938; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_79 = _T_1933[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1940 = $signed(inSpriteY_79) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1941 = _T_1939 & _T_1940; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1942 = $signed(inSpriteY_79) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_80 = $signed(_T_425) - $signed(spriteXPositionReg_80); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1274 = {{1{spriteYPositionReg_80[9]}},spriteYPositionReg_80}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1952 = $signed(_T_431) - $signed(_GEN_1274); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1956 = $signed(inSpriteX_80) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1957 = $signed(inSpriteX_80) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1958 = _T_1956 & _T_1957; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_80 = _T_1952[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1959 = $signed(inSpriteY_80) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1960 = _T_1958 & _T_1959; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1961 = $signed(inSpriteY_80) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_81 = $signed(_T_425) - $signed(spriteXPositionReg_81); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1276 = {{1{spriteYPositionReg_81[9]}},spriteYPositionReg_81}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1971 = $signed(_T_431) - $signed(_GEN_1276); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1975 = $signed(inSpriteX_81) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1976 = $signed(inSpriteX_81) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1977 = _T_1975 & _T_1976; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_81 = _T_1971[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1978 = $signed(inSpriteY_81) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1979 = _T_1977 & _T_1978; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1980 = $signed(inSpriteY_81) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_82 = $signed(_T_425) - $signed(spriteXPositionReg_82); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1278 = {{1{spriteYPositionReg_82[9]}},spriteYPositionReg_82}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_1990 = $signed(_T_431) - $signed(_GEN_1278); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_1994 = $signed(inSpriteX_82) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_1995 = $signed(inSpriteX_82) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_1996 = _T_1994 & _T_1995; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_82 = _T_1990[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_1997 = $signed(inSpriteY_82) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_1998 = _T_1996 & _T_1997; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_1999 = $signed(inSpriteY_82) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_83 = $signed(_T_425) - $signed(spriteXPositionReg_83); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1280 = {{1{spriteYPositionReg_83[9]}},spriteYPositionReg_83}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2009 = $signed(_T_431) - $signed(_GEN_1280); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2013 = $signed(inSpriteX_83) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2014 = $signed(inSpriteX_83) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2015 = _T_2013 & _T_2014; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_83 = _T_2009[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2016 = $signed(inSpriteY_83) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2017 = _T_2015 & _T_2016; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2018 = $signed(inSpriteY_83) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_84 = $signed(_T_425) - $signed(spriteXPositionReg_84); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1282 = {{1{spriteYPositionReg_84[9]}},spriteYPositionReg_84}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2028 = $signed(_T_431) - $signed(_GEN_1282); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2032 = $signed(inSpriteX_84) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2033 = $signed(inSpriteX_84) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2034 = _T_2032 & _T_2033; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_84 = _T_2028[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2035 = $signed(inSpriteY_84) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2036 = _T_2034 & _T_2035; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2037 = $signed(inSpriteY_84) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_85 = $signed(_T_425) - $signed(spriteXPositionReg_85); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1284 = {{1{spriteYPositionReg_85[9]}},spriteYPositionReg_85}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2047 = $signed(_T_431) - $signed(_GEN_1284); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2051 = $signed(inSpriteX_85) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2052 = $signed(inSpriteX_85) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2053 = _T_2051 & _T_2052; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_85 = _T_2047[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2054 = $signed(inSpriteY_85) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2055 = _T_2053 & _T_2054; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2056 = $signed(inSpriteY_85) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_86 = $signed(_T_425) - $signed(spriteXPositionReg_86); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1286 = {{1{spriteYPositionReg_86[9]}},spriteYPositionReg_86}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2066 = $signed(_T_431) - $signed(_GEN_1286); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2070 = $signed(inSpriteX_86) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2071 = $signed(inSpriteX_86) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2072 = _T_2070 & _T_2071; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_86 = _T_2066[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2073 = $signed(inSpriteY_86) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2074 = _T_2072 & _T_2073; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2075 = $signed(inSpriteY_86) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_87 = $signed(_T_425) - $signed(spriteXPositionReg_87); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1288 = {{1{spriteYPositionReg_87[9]}},spriteYPositionReg_87}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2085 = $signed(_T_431) - $signed(_GEN_1288); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2089 = $signed(inSpriteX_87) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2090 = $signed(inSpriteX_87) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2091 = _T_2089 & _T_2090; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_87 = _T_2085[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2092 = $signed(inSpriteY_87) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2093 = _T_2091 & _T_2092; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2094 = $signed(inSpriteY_87) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_88 = $signed(_T_425) - $signed(spriteXPositionReg_88); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1290 = {{1{spriteYPositionReg_88[9]}},spriteYPositionReg_88}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2104 = $signed(_T_431) - $signed(_GEN_1290); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2108 = $signed(inSpriteX_88) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2109 = $signed(inSpriteX_88) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2110 = _T_2108 & _T_2109; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_88 = _T_2104[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2111 = $signed(inSpriteY_88) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2112 = _T_2110 & _T_2111; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2113 = $signed(inSpriteY_88) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_89 = $signed(_T_425) - $signed(spriteXPositionReg_89); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1292 = {{1{spriteYPositionReg_89[9]}},spriteYPositionReg_89}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2123 = $signed(_T_431) - $signed(_GEN_1292); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2127 = $signed(inSpriteX_89) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2128 = $signed(inSpriteX_89) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2129 = _T_2127 & _T_2128; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_89 = _T_2123[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2130 = $signed(inSpriteY_89) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2131 = _T_2129 & _T_2130; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2132 = $signed(inSpriteY_89) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_90 = $signed(_T_425) - $signed(spriteXPositionReg_90); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1294 = {{1{spriteYPositionReg_90[9]}},spriteYPositionReg_90}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2142 = $signed(_T_431) - $signed(_GEN_1294); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2146 = $signed(inSpriteX_90) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2147 = $signed(inSpriteX_90) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2148 = _T_2146 & _T_2147; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_90 = _T_2142[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2149 = $signed(inSpriteY_90) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2150 = _T_2148 & _T_2149; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2151 = $signed(inSpriteY_90) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_91 = $signed(_T_425) - $signed(spriteXPositionReg_91); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1296 = {{1{spriteYPositionReg_91[9]}},spriteYPositionReg_91}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2161 = $signed(_T_431) - $signed(_GEN_1296); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2165 = $signed(inSpriteX_91) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2166 = $signed(inSpriteX_91) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2167 = _T_2165 & _T_2166; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_91 = _T_2161[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2168 = $signed(inSpriteY_91) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2169 = _T_2167 & _T_2168; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2170 = $signed(inSpriteY_91) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_92 = $signed(_T_425) - $signed(spriteXPositionReg_92); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1298 = {{1{spriteYPositionReg_92[9]}},spriteYPositionReg_92}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2180 = $signed(_T_431) - $signed(_GEN_1298); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2184 = $signed(inSpriteX_92) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2185 = $signed(inSpriteX_92) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2186 = _T_2184 & _T_2185; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_92 = _T_2180[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2187 = $signed(inSpriteY_92) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2188 = _T_2186 & _T_2187; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2189 = $signed(inSpriteY_92) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_93 = $signed(_T_425) - $signed(spriteXPositionReg_93); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1300 = {{1{spriteYPositionReg_93[9]}},spriteYPositionReg_93}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2199 = $signed(_T_431) - $signed(_GEN_1300); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2203 = $signed(inSpriteX_93) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2204 = $signed(inSpriteX_93) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2205 = _T_2203 & _T_2204; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_93 = _T_2199[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2206 = $signed(inSpriteY_93) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2207 = _T_2205 & _T_2206; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2208 = $signed(inSpriteY_93) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_94 = $signed(_T_425) - $signed(spriteXPositionReg_94); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1302 = {{1{spriteYPositionReg_94[9]}},spriteYPositionReg_94}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2218 = $signed(_T_431) - $signed(_GEN_1302); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2222 = $signed(inSpriteX_94) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2223 = $signed(inSpriteX_94) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2224 = _T_2222 & _T_2223; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_94 = _T_2218[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2225 = $signed(inSpriteY_94) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2226 = _T_2224 & _T_2225; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2227 = $signed(inSpriteY_94) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_95 = $signed(_T_425) - $signed(spriteXPositionReg_95); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1304 = {{1{spriteYPositionReg_95[9]}},spriteYPositionReg_95}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2237 = $signed(_T_431) - $signed(_GEN_1304); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2241 = $signed(inSpriteX_95) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2242 = $signed(inSpriteX_95) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2243 = _T_2241 & _T_2242; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_95 = _T_2237[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2244 = $signed(inSpriteY_95) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2245 = _T_2243 & _T_2244; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2246 = $signed(inSpriteY_95) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_96 = $signed(_T_425) - $signed(spriteXPositionReg_96); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1306 = {{1{spriteYPositionReg_96[9]}},spriteYPositionReg_96}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2256 = $signed(_T_431) - $signed(_GEN_1306); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2260 = $signed(inSpriteX_96) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2261 = $signed(inSpriteX_96) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2262 = _T_2260 & _T_2261; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_96 = _T_2256[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2263 = $signed(inSpriteY_96) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2264 = _T_2262 & _T_2263; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2265 = $signed(inSpriteY_96) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_97 = $signed(_T_425) - $signed(spriteXPositionReg_97); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1308 = {{1{spriteYPositionReg_97[9]}},spriteYPositionReg_97}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2275 = $signed(_T_431) - $signed(_GEN_1308); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2279 = $signed(inSpriteX_97) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2280 = $signed(inSpriteX_97) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2281 = _T_2279 & _T_2280; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_97 = _T_2275[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2282 = $signed(inSpriteY_97) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2283 = _T_2281 & _T_2282; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2284 = $signed(inSpriteY_97) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_98 = $signed(_T_425) - $signed(spriteXPositionReg_98); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1310 = {{1{spriteYPositionReg_98[9]}},spriteYPositionReg_98}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2294 = $signed(_T_431) - $signed(_GEN_1310); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2298 = $signed(inSpriteX_98) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2299 = $signed(inSpriteX_98) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2300 = _T_2298 & _T_2299; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_98 = _T_2294[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2301 = $signed(inSpriteY_98) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2302 = _T_2300 & _T_2301; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2303 = $signed(inSpriteY_98) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_99 = $signed(_T_425) - $signed(spriteXPositionReg_99); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1312 = {{1{spriteYPositionReg_99[9]}},spriteYPositionReg_99}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2313 = $signed(_T_431) - $signed(_GEN_1312); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2317 = $signed(inSpriteX_99) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2318 = $signed(inSpriteX_99) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2319 = _T_2317 & _T_2318; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_99 = _T_2313[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2320 = $signed(inSpriteY_99) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2321 = _T_2319 & _T_2320; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2322 = $signed(inSpriteY_99) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_100 = $signed(_T_425) - $signed(spriteXPositionReg_100); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1314 = {{1{spriteYPositionReg_100[9]}},spriteYPositionReg_100}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2332 = $signed(_T_431) - $signed(_GEN_1314); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2336 = $signed(inSpriteX_100) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2337 = $signed(inSpriteX_100) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2338 = _T_2336 & _T_2337; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_100 = _T_2332[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2339 = $signed(inSpriteY_100) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2340 = _T_2338 & _T_2339; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2341 = $signed(inSpriteY_100) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_101 = $signed(_T_425) - $signed(spriteXPositionReg_101); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1316 = {{1{spriteYPositionReg_101[9]}},spriteYPositionReg_101}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2351 = $signed(_T_431) - $signed(_GEN_1316); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2355 = $signed(inSpriteX_101) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2356 = $signed(inSpriteX_101) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2357 = _T_2355 & _T_2356; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_101 = _T_2351[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2358 = $signed(inSpriteY_101) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2359 = _T_2357 & _T_2358; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2360 = $signed(inSpriteY_101) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_102 = $signed(_T_425) - $signed(spriteXPositionReg_102); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1318 = {{1{spriteYPositionReg_102[9]}},spriteYPositionReg_102}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2370 = $signed(_T_431) - $signed(_GEN_1318); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2374 = $signed(inSpriteX_102) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2375 = $signed(inSpriteX_102) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2376 = _T_2374 & _T_2375; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_102 = _T_2370[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2377 = $signed(inSpriteY_102) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2378 = _T_2376 & _T_2377; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2379 = $signed(inSpriteY_102) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_103 = $signed(_T_425) - $signed(spriteXPositionReg_103); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1320 = {{1{spriteYPositionReg_103[9]}},spriteYPositionReg_103}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2389 = $signed(_T_431) - $signed(_GEN_1320); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2393 = $signed(inSpriteX_103) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2394 = $signed(inSpriteX_103) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2395 = _T_2393 & _T_2394; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_103 = _T_2389[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2396 = $signed(inSpriteY_103) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2397 = _T_2395 & _T_2396; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2398 = $signed(inSpriteY_103) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_104 = $signed(_T_425) - $signed(spriteXPositionReg_104); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1322 = {{1{spriteYPositionReg_104[9]}},spriteYPositionReg_104}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2408 = $signed(_T_431) - $signed(_GEN_1322); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2412 = $signed(inSpriteX_104) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2413 = $signed(inSpriteX_104) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2414 = _T_2412 & _T_2413; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_104 = _T_2408[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2415 = $signed(inSpriteY_104) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2416 = _T_2414 & _T_2415; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2417 = $signed(inSpriteY_104) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_105 = $signed(_T_425) - $signed(spriteXPositionReg_105); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1324 = {{1{spriteYPositionReg_105[9]}},spriteYPositionReg_105}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2427 = $signed(_T_431) - $signed(_GEN_1324); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2431 = $signed(inSpriteX_105) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2432 = $signed(inSpriteX_105) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2433 = _T_2431 & _T_2432; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_105 = _T_2427[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2434 = $signed(inSpriteY_105) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2435 = _T_2433 & _T_2434; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2436 = $signed(inSpriteY_105) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_106 = $signed(_T_425) - $signed(spriteXPositionReg_106); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1326 = {{1{spriteYPositionReg_106[9]}},spriteYPositionReg_106}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2446 = $signed(_T_431) - $signed(_GEN_1326); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2450 = $signed(inSpriteX_106) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2451 = $signed(inSpriteX_106) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2452 = _T_2450 & _T_2451; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_106 = _T_2446[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2453 = $signed(inSpriteY_106) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2454 = _T_2452 & _T_2453; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2455 = $signed(inSpriteY_106) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_107 = $signed(_T_425) - $signed(spriteXPositionReg_107); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1328 = {{1{spriteYPositionReg_107[9]}},spriteYPositionReg_107}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2465 = $signed(_T_431) - $signed(_GEN_1328); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2469 = $signed(inSpriteX_107) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2470 = $signed(inSpriteX_107) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2471 = _T_2469 & _T_2470; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_107 = _T_2465[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2472 = $signed(inSpriteY_107) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2473 = _T_2471 & _T_2472; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2474 = $signed(inSpriteY_107) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_108 = $signed(_T_425) - $signed(spriteXPositionReg_108); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1330 = {{1{spriteYPositionReg_108[9]}},spriteYPositionReg_108}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2484 = $signed(_T_431) - $signed(_GEN_1330); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2488 = $signed(inSpriteX_108) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2489 = $signed(inSpriteX_108) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2490 = _T_2488 & _T_2489; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_108 = _T_2484[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2491 = $signed(inSpriteY_108) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2492 = _T_2490 & _T_2491; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2493 = $signed(inSpriteY_108) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_109 = $signed(_T_425) - $signed(spriteXPositionReg_109); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1332 = {{1{spriteYPositionReg_109[9]}},spriteYPositionReg_109}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2503 = $signed(_T_431) - $signed(_GEN_1332); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2507 = $signed(inSpriteX_109) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2508 = $signed(inSpriteX_109) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2509 = _T_2507 & _T_2508; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_109 = _T_2503[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2510 = $signed(inSpriteY_109) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2511 = _T_2509 & _T_2510; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2512 = $signed(inSpriteY_109) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_110 = $signed(_T_425) - $signed(spriteXPositionReg_110); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1334 = {{1{spriteYPositionReg_110[9]}},spriteYPositionReg_110}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2522 = $signed(_T_431) - $signed(_GEN_1334); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2526 = $signed(inSpriteX_110) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2527 = $signed(inSpriteX_110) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2528 = _T_2526 & _T_2527; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_110 = _T_2522[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2529 = $signed(inSpriteY_110) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2530 = _T_2528 & _T_2529; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2531 = $signed(inSpriteY_110) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_111 = $signed(_T_425) - $signed(spriteXPositionReg_111); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1336 = {{1{spriteYPositionReg_111[9]}},spriteYPositionReg_111}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2541 = $signed(_T_431) - $signed(_GEN_1336); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2545 = $signed(inSpriteX_111) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2546 = $signed(inSpriteX_111) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2547 = _T_2545 & _T_2546; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_111 = _T_2541[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2548 = $signed(inSpriteY_111) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2549 = _T_2547 & _T_2548; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2550 = $signed(inSpriteY_111) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_112 = $signed(_T_425) - $signed(spriteXPositionReg_112); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1338 = {{1{spriteYPositionReg_112[9]}},spriteYPositionReg_112}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2560 = $signed(_T_431) - $signed(_GEN_1338); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2564 = $signed(inSpriteX_112) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2565 = $signed(inSpriteX_112) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2566 = _T_2564 & _T_2565; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_112 = _T_2560[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2567 = $signed(inSpriteY_112) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2568 = _T_2566 & _T_2567; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2569 = $signed(inSpriteY_112) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_113 = $signed(_T_425) - $signed(spriteXPositionReg_113); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1340 = {{1{spriteYPositionReg_113[9]}},spriteYPositionReg_113}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2579 = $signed(_T_431) - $signed(_GEN_1340); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2583 = $signed(inSpriteX_113) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2584 = $signed(inSpriteX_113) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2585 = _T_2583 & _T_2584; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_113 = _T_2579[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2586 = $signed(inSpriteY_113) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2587 = _T_2585 & _T_2586; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2588 = $signed(inSpriteY_113) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_114 = $signed(_T_425) - $signed(spriteXPositionReg_114); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1342 = {{1{spriteYPositionReg_114[9]}},spriteYPositionReg_114}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2598 = $signed(_T_431) - $signed(_GEN_1342); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2602 = $signed(inSpriteX_114) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2603 = $signed(inSpriteX_114) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2604 = _T_2602 & _T_2603; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_114 = _T_2598[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2605 = $signed(inSpriteY_114) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2606 = _T_2604 & _T_2605; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2607 = $signed(inSpriteY_114) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_115 = $signed(_T_425) - $signed(spriteXPositionReg_115); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1344 = {{1{spriteYPositionReg_115[9]}},spriteYPositionReg_115}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2617 = $signed(_T_431) - $signed(_GEN_1344); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2621 = $signed(inSpriteX_115) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2622 = $signed(inSpriteX_115) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2623 = _T_2621 & _T_2622; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_115 = _T_2617[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2624 = $signed(inSpriteY_115) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2625 = _T_2623 & _T_2624; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2626 = $signed(inSpriteY_115) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_116 = $signed(_T_425) - $signed(spriteXPositionReg_116); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1346 = {{1{spriteYPositionReg_116[9]}},spriteYPositionReg_116}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2636 = $signed(_T_431) - $signed(_GEN_1346); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2640 = $signed(inSpriteX_116) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2641 = $signed(inSpriteX_116) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2642 = _T_2640 & _T_2641; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_116 = _T_2636[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2643 = $signed(inSpriteY_116) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2644 = _T_2642 & _T_2643; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2645 = $signed(inSpriteY_116) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_117 = $signed(_T_425) - $signed(spriteXPositionReg_117); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1348 = {{1{spriteYPositionReg_117[9]}},spriteYPositionReg_117}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2655 = $signed(_T_431) - $signed(_GEN_1348); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2659 = $signed(inSpriteX_117) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2660 = $signed(inSpriteX_117) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2661 = _T_2659 & _T_2660; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_117 = _T_2655[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2662 = $signed(inSpriteY_117) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2663 = _T_2661 & _T_2662; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2664 = $signed(inSpriteY_117) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_118 = $signed(_T_425) - $signed(spriteXPositionReg_118); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1350 = {{1{spriteYPositionReg_118[9]}},spriteYPositionReg_118}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2674 = $signed(_T_431) - $signed(_GEN_1350); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2678 = $signed(inSpriteX_118) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2679 = $signed(inSpriteX_118) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2680 = _T_2678 & _T_2679; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_118 = _T_2674[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2681 = $signed(inSpriteY_118) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2682 = _T_2680 & _T_2681; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2683 = $signed(inSpriteY_118) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_119 = $signed(_T_425) - $signed(spriteXPositionReg_119); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1352 = {{1{spriteYPositionReg_119[9]}},spriteYPositionReg_119}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2693 = $signed(_T_431) - $signed(_GEN_1352); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2697 = $signed(inSpriteX_119) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2698 = $signed(inSpriteX_119) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2699 = _T_2697 & _T_2698; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_119 = _T_2693[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2700 = $signed(inSpriteY_119) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2701 = _T_2699 & _T_2700; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2702 = $signed(inSpriteY_119) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_120 = $signed(_T_425) - $signed(spriteXPositionReg_120); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1354 = {{1{spriteYPositionReg_120[9]}},spriteYPositionReg_120}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2712 = $signed(_T_431) - $signed(_GEN_1354); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2716 = $signed(inSpriteX_120) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2717 = $signed(inSpriteX_120) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2718 = _T_2716 & _T_2717; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_120 = _T_2712[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2719 = $signed(inSpriteY_120) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2720 = _T_2718 & _T_2719; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2721 = $signed(inSpriteY_120) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_121 = $signed(_T_425) - $signed(spriteXPositionReg_121); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1356 = {{1{spriteYPositionReg_121[9]}},spriteYPositionReg_121}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2731 = $signed(_T_431) - $signed(_GEN_1356); // @[GraphicEngineVGA.scala 287:54]
  wire  _T_2735 = $signed(inSpriteX_121) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2736 = $signed(inSpriteX_121) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2737 = _T_2735 & _T_2736; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_121 = _T_2731[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2738 = $signed(inSpriteY_121) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2739 = _T_2737 & _T_2738; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2740 = $signed(inSpriteY_121) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_122 = $signed(_T_425) - $signed(spriteXPositionReg_122); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1358 = {{1{spriteYPositionReg_122[9]}},spriteYPositionReg_122}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2750 = $signed(_T_431) - $signed(_GEN_1358); // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2753 = 12'sh1f - $signed(_T_2750); // @[GraphicEngineVGA.scala 289:28]
  wire [11:0] _GEN_979 = spriteFlipVerticalReg_122 ? $signed(_T_2753) : $signed(_T_2750); // @[GraphicEngineVGA.scala 288:35]
  wire  _T_2754 = $signed(inSpriteX_122) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2755 = $signed(inSpriteX_122) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2756 = _T_2754 & _T_2755; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_122 = _GEN_979[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2757 = $signed(inSpriteY_122) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2758 = _T_2756 & _T_2757; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2759 = $signed(inSpriteY_122) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_123 = $signed(_T_425) - $signed(spriteXPositionReg_123); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1360 = {{1{spriteYPositionReg_123[9]}},spriteYPositionReg_123}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2769 = $signed(_T_431) - $signed(_GEN_1360); // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2772 = 12'sh1f - $signed(_T_2769); // @[GraphicEngineVGA.scala 289:28]
  wire [11:0] _GEN_981 = spriteFlipVerticalReg_123 ? $signed(_T_2772) : $signed(_T_2769); // @[GraphicEngineVGA.scala 288:35]
  wire  _T_2773 = $signed(inSpriteX_123) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2774 = $signed(inSpriteX_123) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2775 = _T_2773 & _T_2774; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_123 = _GEN_981[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2776 = $signed(inSpriteY_123) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2777 = _T_2775 & _T_2776; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2778 = $signed(inSpriteY_123) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_124 = $signed(_T_425) - $signed(spriteXPositionReg_124); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1362 = {{1{spriteYPositionReg_124[9]}},spriteYPositionReg_124}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2788 = $signed(_T_431) - $signed(_GEN_1362); // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2791 = 12'sh1f - $signed(_T_2788); // @[GraphicEngineVGA.scala 289:28]
  wire [11:0] _GEN_983 = spriteFlipVerticalReg_124 ? $signed(_T_2791) : $signed(_T_2788); // @[GraphicEngineVGA.scala 288:35]
  wire  _T_2792 = $signed(inSpriteX_124) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2793 = $signed(inSpriteX_124) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2794 = _T_2792 & _T_2793; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_124 = _GEN_983[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2795 = $signed(inSpriteY_124) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2796 = _T_2794 & _T_2795; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2797 = $signed(inSpriteY_124) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_125 = $signed(_T_425) - $signed(spriteXPositionReg_125); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1364 = {{1{spriteYPositionReg_125[9]}},spriteYPositionReg_125}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2807 = $signed(_T_431) - $signed(_GEN_1364); // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2810 = 12'sh1f - $signed(_T_2807); // @[GraphicEngineVGA.scala 289:28]
  wire [11:0] _GEN_985 = spriteFlipVerticalReg_125 ? $signed(_T_2810) : $signed(_T_2807); // @[GraphicEngineVGA.scala 288:35]
  wire  _T_2811 = $signed(inSpriteX_125) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2812 = $signed(inSpriteX_125) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2813 = _T_2811 & _T_2812; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_125 = _GEN_985[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2814 = $signed(inSpriteY_125) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2815 = _T_2813 & _T_2814; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2816 = $signed(inSpriteY_125) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_126 = $signed(_T_425) - $signed(spriteXPositionReg_126); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1366 = {{1{spriteYPositionReg_126[9]}},spriteYPositionReg_126}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2826 = $signed(_T_431) - $signed(_GEN_1366); // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2829 = 12'sh1f - $signed(_T_2826); // @[GraphicEngineVGA.scala 289:28]
  wire [11:0] _GEN_987 = spriteFlipVerticalReg_126 ? $signed(_T_2829) : $signed(_T_2826); // @[GraphicEngineVGA.scala 288:35]
  wire  _T_2830 = $signed(inSpriteX_126) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2831 = $signed(inSpriteX_126) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2832 = _T_2830 & _T_2831; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_126 = _GEN_987[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2833 = $signed(inSpriteY_126) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2834 = _T_2832 & _T_2833; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2835 = $signed(inSpriteY_126) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [11:0] inSpriteX_127 = $signed(_T_425) - $signed(spriteXPositionReg_127); // @[GraphicEngineVGA.scala 281:54]
  wire [10:0] _GEN_1368 = {{1{spriteYPositionReg_127[9]}},spriteYPositionReg_127}; // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2845 = $signed(_T_431) - $signed(_GEN_1368); // @[GraphicEngineVGA.scala 287:54]
  wire [11:0] _T_2848 = 12'sh1f - $signed(_T_2845); // @[GraphicEngineVGA.scala 289:28]
  wire [11:0] _GEN_989 = spriteFlipVerticalReg_127 ? $signed(_T_2848) : $signed(_T_2845); // @[GraphicEngineVGA.scala 288:35]
  wire  _T_2849 = $signed(inSpriteX_127) >= 12'sh0; // @[GraphicEngineVGA.scala 293:33]
  wire  _T_2850 = $signed(inSpriteX_127) < 12'sh20; // @[GraphicEngineVGA.scala 293:56]
  wire  _T_2851 = _T_2849 & _T_2850; // @[GraphicEngineVGA.scala 293:40]
  wire [10:0] inSpriteY_127 = _GEN_989[10:0]; // @[GraphicEngineVGA.scala 279:23 GraphicEngineVGA.scala 289:20 GraphicEngineVGA.scala 291:20]
  wire  _T_2852 = $signed(inSpriteY_127) >= 11'sh0; // @[GraphicEngineVGA.scala 293:79]
  wire  _T_2853 = _T_2851 & _T_2852; // @[GraphicEngineVGA.scala 293:63]
  wire  _T_2854 = $signed(inSpriteY_127) < 11'sh20; // @[GraphicEngineVGA.scala 293:102]
  wire [5:0] _GEN_1370 = {{1'd0}, inSpriteY_0[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2858 = 6'h20 * _GEN_1370; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1371 = {{6'd0}, inSpriteX_0[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2860 = _GEN_1371 + _T_2858; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1372 = {{1'd0}, inSpriteY_1[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2863 = 6'h20 * _GEN_1372; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1373 = {{6'd0}, inSpriteX_1[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2865 = _GEN_1373 + _T_2863; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1374 = {{1'd0}, inSpriteY_2[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2868 = 6'h20 * _GEN_1374; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1375 = {{6'd0}, inSpriteX_2[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2870 = _GEN_1375 + _T_2868; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1376 = {{1'd0}, inSpriteY_3[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2873 = 6'h20 * _GEN_1376; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1377 = {{6'd0}, inSpriteX_3[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2875 = _GEN_1377 + _T_2873; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1378 = {{1'd0}, inSpriteY_4[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2878 = 6'h20 * _GEN_1378; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1379 = {{6'd0}, inSpriteX_4[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2880 = _GEN_1379 + _T_2878; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1380 = {{1'd0}, inSpriteY_5[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2883 = 6'h20 * _GEN_1380; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1381 = {{6'd0}, inSpriteX_5[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2885 = _GEN_1381 + _T_2883; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1382 = {{1'd0}, inSpriteY_6[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2888 = 6'h20 * _GEN_1382; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1383 = {{6'd0}, inSpriteX_6[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2890 = _GEN_1383 + _T_2888; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1384 = {{1'd0}, inSpriteY_7[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2893 = 6'h20 * _GEN_1384; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1385 = {{6'd0}, inSpriteX_7[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2895 = _GEN_1385 + _T_2893; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1386 = {{1'd0}, inSpriteY_8[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2898 = 6'h20 * _GEN_1386; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1387 = {{6'd0}, inSpriteX_8[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2900 = _GEN_1387 + _T_2898; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1388 = {{1'd0}, inSpriteY_9[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2903 = 6'h20 * _GEN_1388; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1389 = {{6'd0}, inSpriteX_9[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2905 = _GEN_1389 + _T_2903; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1390 = {{1'd0}, inSpriteY_10[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2908 = 6'h20 * _GEN_1390; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1391 = {{6'd0}, inSpriteX_10[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2910 = _GEN_1391 + _T_2908; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1392 = {{1'd0}, inSpriteY_11[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2913 = 6'h20 * _GEN_1392; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1393 = {{6'd0}, inSpriteX_11[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2915 = _GEN_1393 + _T_2913; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1394 = {{1'd0}, inSpriteY_12[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2918 = 6'h20 * _GEN_1394; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1395 = {{6'd0}, inSpriteX_12[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2920 = _GEN_1395 + _T_2918; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1396 = {{1'd0}, inSpriteY_13[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2923 = 6'h20 * _GEN_1396; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1397 = {{6'd0}, inSpriteX_13[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2925 = _GEN_1397 + _T_2923; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1398 = {{1'd0}, inSpriteY_14[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2928 = 6'h20 * _GEN_1398; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1399 = {{6'd0}, inSpriteX_14[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2930 = _GEN_1399 + _T_2928; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1400 = {{1'd0}, inSpriteY_15[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2933 = 6'h20 * _GEN_1400; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1401 = {{6'd0}, inSpriteX_15[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2935 = _GEN_1401 + _T_2933; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1402 = {{1'd0}, inSpriteY_16[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2938 = 6'h20 * _GEN_1402; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1403 = {{6'd0}, inSpriteX_16[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2940 = _GEN_1403 + _T_2938; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1404 = {{1'd0}, inSpriteY_17[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2943 = 6'h20 * _GEN_1404; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1405 = {{6'd0}, inSpriteX_17[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2945 = _GEN_1405 + _T_2943; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1406 = {{1'd0}, inSpriteY_18[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2948 = 6'h20 * _GEN_1406; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1407 = {{6'd0}, inSpriteX_18[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2950 = _GEN_1407 + _T_2948; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1408 = {{1'd0}, inSpriteY_19[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2953 = 6'h20 * _GEN_1408; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1409 = {{6'd0}, inSpriteX_19[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2955 = _GEN_1409 + _T_2953; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1410 = {{1'd0}, inSpriteY_20[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2958 = 6'h20 * _GEN_1410; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1411 = {{6'd0}, inSpriteX_20[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2960 = _GEN_1411 + _T_2958; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1412 = {{1'd0}, inSpriteY_21[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2963 = 6'h20 * _GEN_1412; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1413 = {{6'd0}, inSpriteX_21[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2965 = _GEN_1413 + _T_2963; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1414 = {{1'd0}, inSpriteY_22[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2968 = 6'h20 * _GEN_1414; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1415 = {{6'd0}, inSpriteX_22[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2970 = _GEN_1415 + _T_2968; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1416 = {{1'd0}, inSpriteY_23[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2973 = 6'h20 * _GEN_1416; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1417 = {{6'd0}, inSpriteX_23[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2975 = _GEN_1417 + _T_2973; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1418 = {{1'd0}, inSpriteY_24[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2978 = 6'h20 * _GEN_1418; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1419 = {{6'd0}, inSpriteX_24[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2980 = _GEN_1419 + _T_2978; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1420 = {{1'd0}, inSpriteY_25[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2983 = 6'h20 * _GEN_1420; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1421 = {{6'd0}, inSpriteX_25[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2985 = _GEN_1421 + _T_2983; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1422 = {{1'd0}, inSpriteY_26[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2988 = 6'h20 * _GEN_1422; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1423 = {{6'd0}, inSpriteX_26[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2990 = _GEN_1423 + _T_2988; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1424 = {{1'd0}, inSpriteY_27[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2993 = 6'h20 * _GEN_1424; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1425 = {{6'd0}, inSpriteX_27[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_2995 = _GEN_1425 + _T_2993; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1426 = {{1'd0}, inSpriteY_28[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_2998 = 6'h20 * _GEN_1426; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1427 = {{6'd0}, inSpriteX_28[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3000 = _GEN_1427 + _T_2998; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1428 = {{1'd0}, inSpriteY_29[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3003 = 6'h20 * _GEN_1428; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1429 = {{6'd0}, inSpriteX_29[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3005 = _GEN_1429 + _T_3003; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1430 = {{1'd0}, inSpriteY_30[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3008 = 6'h20 * _GEN_1430; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1431 = {{6'd0}, inSpriteX_30[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3010 = _GEN_1431 + _T_3008; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1432 = {{1'd0}, inSpriteY_31[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3013 = 6'h20 * _GEN_1432; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1433 = {{6'd0}, inSpriteX_31[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3015 = _GEN_1433 + _T_3013; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1434 = {{1'd0}, inSpriteY_32[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3018 = 6'h20 * _GEN_1434; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1435 = {{6'd0}, inSpriteX_32[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3020 = _GEN_1435 + _T_3018; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1436 = {{1'd0}, inSpriteY_33[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3023 = 6'h20 * _GEN_1436; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1437 = {{6'd0}, inSpriteX_33[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3025 = _GEN_1437 + _T_3023; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1438 = {{1'd0}, inSpriteY_34[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3028 = 6'h20 * _GEN_1438; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1439 = {{6'd0}, inSpriteX_34[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3030 = _GEN_1439 + _T_3028; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1440 = {{1'd0}, inSpriteY_35[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3033 = 6'h20 * _GEN_1440; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1441 = {{6'd0}, inSpriteX_35[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3035 = _GEN_1441 + _T_3033; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1442 = {{1'd0}, inSpriteY_36[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3038 = 6'h20 * _GEN_1442; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1443 = {{6'd0}, inSpriteX_36[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3040 = _GEN_1443 + _T_3038; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1444 = {{1'd0}, inSpriteY_37[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3043 = 6'h20 * _GEN_1444; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1445 = {{6'd0}, inSpriteX_37[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3045 = _GEN_1445 + _T_3043; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1446 = {{1'd0}, inSpriteY_38[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3048 = 6'h20 * _GEN_1446; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1447 = {{6'd0}, inSpriteX_38[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3050 = _GEN_1447 + _T_3048; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1448 = {{1'd0}, inSpriteY_39[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3053 = 6'h20 * _GEN_1448; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1449 = {{6'd0}, inSpriteX_39[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3055 = _GEN_1449 + _T_3053; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1450 = {{1'd0}, inSpriteY_40[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3058 = 6'h20 * _GEN_1450; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1451 = {{6'd0}, inSpriteX_40[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3060 = _GEN_1451 + _T_3058; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1452 = {{1'd0}, inSpriteY_41[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3063 = 6'h20 * _GEN_1452; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1453 = {{6'd0}, inSpriteX_41[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3065 = _GEN_1453 + _T_3063; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1454 = {{1'd0}, inSpriteY_42[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3068 = 6'h20 * _GEN_1454; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1455 = {{6'd0}, inSpriteX_42[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3070 = _GEN_1455 + _T_3068; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1456 = {{1'd0}, inSpriteY_43[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3073 = 6'h20 * _GEN_1456; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1457 = {{6'd0}, inSpriteX_43[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3075 = _GEN_1457 + _T_3073; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1458 = {{1'd0}, inSpriteY_44[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3078 = 6'h20 * _GEN_1458; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1459 = {{6'd0}, inSpriteX_44[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3080 = _GEN_1459 + _T_3078; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1460 = {{1'd0}, inSpriteY_45[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3083 = 6'h20 * _GEN_1460; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1461 = {{6'd0}, inSpriteX_45[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3085 = _GEN_1461 + _T_3083; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1462 = {{1'd0}, inSpriteY_46[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3088 = 6'h20 * _GEN_1462; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1463 = {{6'd0}, inSpriteX_46[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3090 = _GEN_1463 + _T_3088; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1464 = {{1'd0}, inSpriteY_47[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3093 = 6'h20 * _GEN_1464; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1465 = {{6'd0}, inSpriteX_47[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3095 = _GEN_1465 + _T_3093; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1466 = {{1'd0}, inSpriteY_48[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3098 = 6'h20 * _GEN_1466; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1467 = {{6'd0}, inSpriteX_48[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3100 = _GEN_1467 + _T_3098; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1468 = {{1'd0}, inSpriteY_49[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3103 = 6'h20 * _GEN_1468; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1469 = {{6'd0}, inSpriteX_49[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3105 = _GEN_1469 + _T_3103; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1470 = {{1'd0}, inSpriteY_50[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3108 = 6'h20 * _GEN_1470; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1471 = {{6'd0}, inSpriteX_50[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3110 = _GEN_1471 + _T_3108; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1472 = {{1'd0}, inSpriteY_51[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3113 = 6'h20 * _GEN_1472; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1473 = {{6'd0}, inSpriteX_51[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3115 = _GEN_1473 + _T_3113; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1474 = {{1'd0}, inSpriteY_52[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3118 = 6'h20 * _GEN_1474; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1475 = {{6'd0}, inSpriteX_52[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3120 = _GEN_1475 + _T_3118; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1476 = {{1'd0}, inSpriteY_53[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3123 = 6'h20 * _GEN_1476; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1477 = {{6'd0}, inSpriteX_53[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3125 = _GEN_1477 + _T_3123; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1478 = {{1'd0}, inSpriteY_54[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3128 = 6'h20 * _GEN_1478; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1479 = {{6'd0}, inSpriteX_54[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3130 = _GEN_1479 + _T_3128; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1480 = {{1'd0}, inSpriteY_55[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3133 = 6'h20 * _GEN_1480; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1481 = {{6'd0}, inSpriteX_55[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3135 = _GEN_1481 + _T_3133; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1482 = {{1'd0}, inSpriteY_56[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3138 = 6'h20 * _GEN_1482; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1483 = {{6'd0}, inSpriteX_56[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3140 = _GEN_1483 + _T_3138; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1484 = {{1'd0}, inSpriteY_57[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3143 = 6'h20 * _GEN_1484; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1485 = {{6'd0}, inSpriteX_57[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3145 = _GEN_1485 + _T_3143; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1486 = {{1'd0}, inSpriteY_58[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3148 = 6'h20 * _GEN_1486; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1487 = {{6'd0}, inSpriteX_58[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3150 = _GEN_1487 + _T_3148; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1488 = {{1'd0}, inSpriteY_59[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3153 = 6'h20 * _GEN_1488; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1489 = {{6'd0}, inSpriteX_59[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3155 = _GEN_1489 + _T_3153; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1490 = {{1'd0}, inSpriteY_60[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3158 = 6'h20 * _GEN_1490; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1491 = {{6'd0}, inSpriteX_60[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3160 = _GEN_1491 + _T_3158; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1492 = {{1'd0}, inSpriteY_61[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3163 = 6'h20 * _GEN_1492; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1493 = {{6'd0}, inSpriteX_61[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3165 = _GEN_1493 + _T_3163; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1494 = {{1'd0}, inSpriteY_62[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3168 = 6'h20 * _GEN_1494; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1495 = {{6'd0}, inSpriteX_62[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3170 = _GEN_1495 + _T_3168; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1496 = {{1'd0}, inSpriteY_63[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3173 = 6'h20 * _GEN_1496; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1497 = {{6'd0}, inSpriteX_63[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3175 = _GEN_1497 + _T_3173; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1498 = {{1'd0}, inSpriteY_64[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3178 = 6'h20 * _GEN_1498; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1499 = {{6'd0}, inSpriteX_64[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3180 = _GEN_1499 + _T_3178; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _GEN_1501 = {{6'd0}, inSpriteX_65[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3185 = _GEN_1501 + _T_3178; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _GEN_1503 = {{6'd0}, inSpriteX_66[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3190 = _GEN_1503 + _T_3178; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _GEN_1505 = {{6'd0}, inSpriteX_67[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3195 = _GEN_1505 + _T_3178; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _GEN_1507 = {{6'd0}, inSpriteX_68[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3200 = _GEN_1507 + _T_3178; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _GEN_1509 = {{6'd0}, inSpriteX_69[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3205 = _GEN_1509 + _T_3178; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1510 = {{1'd0}, inSpriteY_70[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3208 = 6'h20 * _GEN_1510; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1511 = {{6'd0}, inSpriteX_70[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3210 = _GEN_1511 + _T_3208; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1512 = {{1'd0}, inSpriteY_71[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3213 = 6'h20 * _GEN_1512; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1513 = {{6'd0}, inSpriteX_71[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3215 = _GEN_1513 + _T_3213; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1514 = {{1'd0}, inSpriteY_72[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3218 = 6'h20 * _GEN_1514; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1515 = {{6'd0}, inSpriteX_72[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3220 = _GEN_1515 + _T_3218; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1516 = {{1'd0}, inSpriteY_73[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3223 = 6'h20 * _GEN_1516; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1517 = {{6'd0}, inSpriteX_73[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3225 = _GEN_1517 + _T_3223; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1518 = {{1'd0}, inSpriteY_74[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3228 = 6'h20 * _GEN_1518; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1519 = {{6'd0}, inSpriteX_74[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3230 = _GEN_1519 + _T_3228; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1520 = {{1'd0}, inSpriteY_75[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3233 = 6'h20 * _GEN_1520; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1521 = {{6'd0}, inSpriteX_75[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3235 = _GEN_1521 + _T_3233; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1522 = {{1'd0}, inSpriteY_76[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3238 = 6'h20 * _GEN_1522; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1523 = {{6'd0}, inSpriteX_76[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3240 = _GEN_1523 + _T_3238; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1524 = {{1'd0}, inSpriteY_77[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3243 = 6'h20 * _GEN_1524; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1525 = {{6'd0}, inSpriteX_77[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3245 = _GEN_1525 + _T_3243; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1526 = {{1'd0}, inSpriteY_78[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3248 = 6'h20 * _GEN_1526; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1527 = {{6'd0}, inSpriteX_78[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3250 = _GEN_1527 + _T_3248; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1528 = {{1'd0}, inSpriteY_79[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3253 = 6'h20 * _GEN_1528; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1529 = {{6'd0}, inSpriteX_79[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3255 = _GEN_1529 + _T_3253; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1530 = {{1'd0}, inSpriteY_80[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3258 = 6'h20 * _GEN_1530; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1531 = {{6'd0}, inSpriteX_80[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3260 = _GEN_1531 + _T_3258; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1532 = {{1'd0}, inSpriteY_81[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3263 = 6'h20 * _GEN_1532; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1533 = {{6'd0}, inSpriteX_81[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3265 = _GEN_1533 + _T_3263; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1534 = {{1'd0}, inSpriteY_82[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3268 = 6'h20 * _GEN_1534; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1535 = {{6'd0}, inSpriteX_82[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3270 = _GEN_1535 + _T_3268; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1536 = {{1'd0}, inSpriteY_83[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3273 = 6'h20 * _GEN_1536; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1537 = {{6'd0}, inSpriteX_83[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3275 = _GEN_1537 + _T_3273; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1538 = {{1'd0}, inSpriteY_84[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3278 = 6'h20 * _GEN_1538; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1539 = {{6'd0}, inSpriteX_84[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3280 = _GEN_1539 + _T_3278; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1540 = {{1'd0}, inSpriteY_85[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3283 = 6'h20 * _GEN_1540; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1541 = {{6'd0}, inSpriteX_85[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3285 = _GEN_1541 + _T_3283; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1542 = {{1'd0}, inSpriteY_86[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3288 = 6'h20 * _GEN_1542; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1543 = {{6'd0}, inSpriteX_86[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3290 = _GEN_1543 + _T_3288; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1544 = {{1'd0}, inSpriteY_87[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3293 = 6'h20 * _GEN_1544; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1545 = {{6'd0}, inSpriteX_87[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3295 = _GEN_1545 + _T_3293; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1546 = {{1'd0}, inSpriteY_88[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3298 = 6'h20 * _GEN_1546; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1547 = {{6'd0}, inSpriteX_88[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3300 = _GEN_1547 + _T_3298; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1548 = {{1'd0}, inSpriteY_89[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3303 = 6'h20 * _GEN_1548; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1549 = {{6'd0}, inSpriteX_89[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3305 = _GEN_1549 + _T_3303; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1550 = {{1'd0}, inSpriteY_90[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3308 = 6'h20 * _GEN_1550; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1551 = {{6'd0}, inSpriteX_90[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3310 = _GEN_1551 + _T_3308; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1552 = {{1'd0}, inSpriteY_91[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3313 = 6'h20 * _GEN_1552; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1553 = {{6'd0}, inSpriteX_91[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3315 = _GEN_1553 + _T_3313; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1554 = {{1'd0}, inSpriteY_92[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3318 = 6'h20 * _GEN_1554; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1555 = {{6'd0}, inSpriteX_92[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3320 = _GEN_1555 + _T_3318; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1556 = {{1'd0}, inSpriteY_93[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3323 = 6'h20 * _GEN_1556; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1557 = {{6'd0}, inSpriteX_93[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3325 = _GEN_1557 + _T_3323; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1558 = {{1'd0}, inSpriteY_94[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3328 = 6'h20 * _GEN_1558; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1559 = {{6'd0}, inSpriteX_94[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3330 = _GEN_1559 + _T_3328; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1560 = {{1'd0}, inSpriteY_95[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3333 = 6'h20 * _GEN_1560; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1561 = {{6'd0}, inSpriteX_95[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3335 = _GEN_1561 + _T_3333; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1562 = {{1'd0}, inSpriteY_96[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3338 = 6'h20 * _GEN_1562; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1563 = {{6'd0}, inSpriteX_96[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3340 = _GEN_1563 + _T_3338; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1564 = {{1'd0}, inSpriteY_97[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3343 = 6'h20 * _GEN_1564; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1565 = {{6'd0}, inSpriteX_97[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3345 = _GEN_1565 + _T_3343; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1566 = {{1'd0}, inSpriteY_98[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3348 = 6'h20 * _GEN_1566; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1567 = {{6'd0}, inSpriteX_98[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3350 = _GEN_1567 + _T_3348; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1568 = {{1'd0}, inSpriteY_99[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3353 = 6'h20 * _GEN_1568; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1569 = {{6'd0}, inSpriteX_99[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3355 = _GEN_1569 + _T_3353; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1570 = {{1'd0}, inSpriteY_100[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3358 = 6'h20 * _GEN_1570; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1571 = {{6'd0}, inSpriteX_100[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3360 = _GEN_1571 + _T_3358; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1572 = {{1'd0}, inSpriteY_101[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3363 = 6'h20 * _GEN_1572; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1573 = {{6'd0}, inSpriteX_101[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3365 = _GEN_1573 + _T_3363; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1574 = {{1'd0}, inSpriteY_102[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3368 = 6'h20 * _GEN_1574; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1575 = {{6'd0}, inSpriteX_102[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3370 = _GEN_1575 + _T_3368; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1576 = {{1'd0}, inSpriteY_103[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3373 = 6'h20 * _GEN_1576; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1577 = {{6'd0}, inSpriteX_103[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3375 = _GEN_1577 + _T_3373; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1578 = {{1'd0}, inSpriteY_104[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3378 = 6'h20 * _GEN_1578; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1579 = {{6'd0}, inSpriteX_104[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3380 = _GEN_1579 + _T_3378; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1580 = {{1'd0}, inSpriteY_105[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3383 = 6'h20 * _GEN_1580; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1581 = {{6'd0}, inSpriteX_105[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3385 = _GEN_1581 + _T_3383; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1582 = {{1'd0}, inSpriteY_106[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3388 = 6'h20 * _GEN_1582; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1583 = {{6'd0}, inSpriteX_106[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3390 = _GEN_1583 + _T_3388; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1584 = {{1'd0}, inSpriteY_107[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3393 = 6'h20 * _GEN_1584; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1585 = {{6'd0}, inSpriteX_107[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3395 = _GEN_1585 + _T_3393; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1586 = {{1'd0}, inSpriteY_108[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3398 = 6'h20 * _GEN_1586; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1587 = {{6'd0}, inSpriteX_108[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3400 = _GEN_1587 + _T_3398; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1588 = {{1'd0}, inSpriteY_109[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3403 = 6'h20 * _GEN_1588; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1589 = {{6'd0}, inSpriteX_109[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3405 = _GEN_1589 + _T_3403; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1590 = {{1'd0}, inSpriteY_110[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3408 = 6'h20 * _GEN_1590; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1591 = {{6'd0}, inSpriteX_110[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3410 = _GEN_1591 + _T_3408; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1592 = {{1'd0}, inSpriteY_111[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3413 = 6'h20 * _GEN_1592; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1593 = {{6'd0}, inSpriteX_111[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3415 = _GEN_1593 + _T_3413; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1594 = {{1'd0}, inSpriteY_112[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3418 = 6'h20 * _GEN_1594; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1595 = {{6'd0}, inSpriteX_112[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3420 = _GEN_1595 + _T_3418; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1596 = {{1'd0}, inSpriteY_113[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3423 = 6'h20 * _GEN_1596; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1597 = {{6'd0}, inSpriteX_113[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3425 = _GEN_1597 + _T_3423; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1598 = {{1'd0}, inSpriteY_114[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3428 = 6'h20 * _GEN_1598; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1599 = {{6'd0}, inSpriteX_114[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3430 = _GEN_1599 + _T_3428; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1600 = {{1'd0}, inSpriteY_115[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3433 = 6'h20 * _GEN_1600; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1601 = {{6'd0}, inSpriteX_115[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3435 = _GEN_1601 + _T_3433; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1602 = {{1'd0}, inSpriteY_116[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3438 = 6'h20 * _GEN_1602; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1603 = {{6'd0}, inSpriteX_116[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3440 = _GEN_1603 + _T_3438; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1604 = {{1'd0}, inSpriteY_117[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3443 = 6'h20 * _GEN_1604; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1605 = {{6'd0}, inSpriteX_117[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3445 = _GEN_1605 + _T_3443; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1606 = {{1'd0}, inSpriteY_118[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3448 = 6'h20 * _GEN_1606; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1607 = {{6'd0}, inSpriteX_118[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3450 = _GEN_1607 + _T_3448; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1608 = {{1'd0}, inSpriteY_119[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3453 = 6'h20 * _GEN_1608; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1609 = {{6'd0}, inSpriteX_119[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3455 = _GEN_1609 + _T_3453; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1610 = {{1'd0}, inSpriteY_120[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3458 = 6'h20 * _GEN_1610; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1611 = {{6'd0}, inSpriteX_120[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3460 = _GEN_1611 + _T_3458; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1612 = {{1'd0}, inSpriteY_121[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3463 = 6'h20 * _GEN_1612; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1613 = {{6'd0}, inSpriteX_121[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3465 = _GEN_1613 + _T_3463; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1614 = {{1'd0}, inSpriteY_122[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3468 = 6'h20 * _GEN_1614; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1615 = {{6'd0}, inSpriteX_122[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3470 = _GEN_1615 + _T_3468; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1616 = {{1'd0}, inSpriteY_123[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3473 = 6'h20 * _GEN_1616; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1617 = {{6'd0}, inSpriteX_123[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3475 = _GEN_1617 + _T_3473; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1618 = {{1'd0}, inSpriteY_124[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3478 = 6'h20 * _GEN_1618; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1619 = {{6'd0}, inSpriteX_124[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3480 = _GEN_1619 + _T_3478; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1620 = {{1'd0}, inSpriteY_125[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3483 = 6'h20 * _GEN_1620; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1621 = {{6'd0}, inSpriteX_125[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3485 = _GEN_1621 + _T_3483; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1622 = {{1'd0}, inSpriteY_126[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3488 = 6'h20 * _GEN_1622; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1623 = {{6'd0}, inSpriteX_126[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3490 = _GEN_1623 + _T_3488; // @[GraphicEngineVGA.scala 301:62]
  wire [5:0] _GEN_1624 = {{1'd0}, inSpriteY_127[4:0]}; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _T_3493 = 6'h20 * _GEN_1624; // @[GraphicEngineVGA.scala 301:74]
  wire [10:0] _GEN_1625 = {{6'd0}, inSpriteX_127[4:0]}; // @[GraphicEngineVGA.scala 301:62]
  wire [10:0] _T_3495 = _GEN_1625 + _T_3493; // @[GraphicEngineVGA.scala 301:62]
  reg [5:0] _T_3497; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3498_0; // @[GameUtilities.scala 21:24]
  reg  _T_3498_1; // @[GameUtilities.scala 21:24]
  reg  _T_3499_0; // @[GameUtilities.scala 21:24]
  reg  _T_3499_1; // @[GameUtilities.scala 21:24]
  wire  _T_3500 = _T_3498_0 & _T_3499_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3502; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3503 = ~_T_3502; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3506; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3507_0; // @[GameUtilities.scala 21:24]
  reg  _T_3507_1; // @[GameUtilities.scala 21:24]
  reg  _T_3508_0; // @[GameUtilities.scala 21:24]
  reg  _T_3508_1; // @[GameUtilities.scala 21:24]
  wire  _T_3509 = _T_3507_0 & _T_3508_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3511; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3512 = ~_T_3511; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3515; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3516_0; // @[GameUtilities.scala 21:24]
  reg  _T_3516_1; // @[GameUtilities.scala 21:24]
  reg  _T_3517_0; // @[GameUtilities.scala 21:24]
  reg  _T_3517_1; // @[GameUtilities.scala 21:24]
  wire  _T_3518 = _T_3516_0 & _T_3517_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3520; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3521 = ~_T_3520; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3524; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3525_0; // @[GameUtilities.scala 21:24]
  reg  _T_3525_1; // @[GameUtilities.scala 21:24]
  reg  _T_3526_0; // @[GameUtilities.scala 21:24]
  reg  _T_3526_1; // @[GameUtilities.scala 21:24]
  wire  _T_3527 = _T_3525_0 & _T_3526_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3529; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3530 = ~_T_3529; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3533; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3534_0; // @[GameUtilities.scala 21:24]
  reg  _T_3534_1; // @[GameUtilities.scala 21:24]
  reg  _T_3535_0; // @[GameUtilities.scala 21:24]
  reg  _T_3535_1; // @[GameUtilities.scala 21:24]
  wire  _T_3536 = _T_3534_0 & _T_3535_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3538; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3539 = ~_T_3538; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3542; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3543_0; // @[GameUtilities.scala 21:24]
  reg  _T_3543_1; // @[GameUtilities.scala 21:24]
  reg  _T_3544_0; // @[GameUtilities.scala 21:24]
  reg  _T_3544_1; // @[GameUtilities.scala 21:24]
  wire  _T_3545 = _T_3543_0 & _T_3544_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3547; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3548 = ~_T_3547; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3551; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3552_0; // @[GameUtilities.scala 21:24]
  reg  _T_3552_1; // @[GameUtilities.scala 21:24]
  reg  _T_3553_0; // @[GameUtilities.scala 21:24]
  reg  _T_3553_1; // @[GameUtilities.scala 21:24]
  wire  _T_3554 = _T_3552_0 & _T_3553_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3556; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3557 = ~_T_3556; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3560; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3561_0; // @[GameUtilities.scala 21:24]
  reg  _T_3561_1; // @[GameUtilities.scala 21:24]
  reg  _T_3562_0; // @[GameUtilities.scala 21:24]
  reg  _T_3562_1; // @[GameUtilities.scala 21:24]
  wire  _T_3563 = _T_3561_0 & _T_3562_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3565; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3566 = ~_T_3565; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3569; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3570_0; // @[GameUtilities.scala 21:24]
  reg  _T_3570_1; // @[GameUtilities.scala 21:24]
  reg  _T_3571_0; // @[GameUtilities.scala 21:24]
  reg  _T_3571_1; // @[GameUtilities.scala 21:24]
  wire  _T_3572 = _T_3570_0 & _T_3571_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3574; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3575 = ~_T_3574; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3578; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3579_0; // @[GameUtilities.scala 21:24]
  reg  _T_3579_1; // @[GameUtilities.scala 21:24]
  reg  _T_3580_0; // @[GameUtilities.scala 21:24]
  reg  _T_3580_1; // @[GameUtilities.scala 21:24]
  wire  _T_3581 = _T_3579_0 & _T_3580_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3583; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3584 = ~_T_3583; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3587; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3588_0; // @[GameUtilities.scala 21:24]
  reg  _T_3588_1; // @[GameUtilities.scala 21:24]
  reg  _T_3589_0; // @[GameUtilities.scala 21:24]
  reg  _T_3589_1; // @[GameUtilities.scala 21:24]
  wire  _T_3590 = _T_3588_0 & _T_3589_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3592; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3593 = ~_T_3592; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3596; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3597_0; // @[GameUtilities.scala 21:24]
  reg  _T_3597_1; // @[GameUtilities.scala 21:24]
  reg  _T_3598_0; // @[GameUtilities.scala 21:24]
  reg  _T_3598_1; // @[GameUtilities.scala 21:24]
  wire  _T_3599 = _T_3597_0 & _T_3598_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3601; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3602 = ~_T_3601; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3605; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3606_0; // @[GameUtilities.scala 21:24]
  reg  _T_3606_1; // @[GameUtilities.scala 21:24]
  reg  _T_3607_0; // @[GameUtilities.scala 21:24]
  reg  _T_3607_1; // @[GameUtilities.scala 21:24]
  wire  _T_3608 = _T_3606_0 & _T_3607_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3610; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3611 = ~_T_3610; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3614; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3615_0; // @[GameUtilities.scala 21:24]
  reg  _T_3615_1; // @[GameUtilities.scala 21:24]
  reg  _T_3616_0; // @[GameUtilities.scala 21:24]
  reg  _T_3616_1; // @[GameUtilities.scala 21:24]
  wire  _T_3617 = _T_3615_0 & _T_3616_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3619; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3620 = ~_T_3619; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3623; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3624_0; // @[GameUtilities.scala 21:24]
  reg  _T_3624_1; // @[GameUtilities.scala 21:24]
  reg  _T_3625_0; // @[GameUtilities.scala 21:24]
  reg  _T_3625_1; // @[GameUtilities.scala 21:24]
  wire  _T_3626 = _T_3624_0 & _T_3625_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3628; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3629 = ~_T_3628; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3632; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3633_0; // @[GameUtilities.scala 21:24]
  reg  _T_3633_1; // @[GameUtilities.scala 21:24]
  reg  _T_3634_0; // @[GameUtilities.scala 21:24]
  reg  _T_3634_1; // @[GameUtilities.scala 21:24]
  wire  _T_3635 = _T_3633_0 & _T_3634_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3637; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3638 = ~_T_3637; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3641; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3642_0; // @[GameUtilities.scala 21:24]
  reg  _T_3642_1; // @[GameUtilities.scala 21:24]
  reg  _T_3643_0; // @[GameUtilities.scala 21:24]
  reg  _T_3643_1; // @[GameUtilities.scala 21:24]
  wire  _T_3644 = _T_3642_0 & _T_3643_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3646; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3647 = ~_T_3646; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3650; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3651_0; // @[GameUtilities.scala 21:24]
  reg  _T_3651_1; // @[GameUtilities.scala 21:24]
  reg  _T_3652_0; // @[GameUtilities.scala 21:24]
  reg  _T_3652_1; // @[GameUtilities.scala 21:24]
  wire  _T_3653 = _T_3651_0 & _T_3652_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3655; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3656 = ~_T_3655; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3659; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3660_0; // @[GameUtilities.scala 21:24]
  reg  _T_3660_1; // @[GameUtilities.scala 21:24]
  reg  _T_3661_0; // @[GameUtilities.scala 21:24]
  reg  _T_3661_1; // @[GameUtilities.scala 21:24]
  wire  _T_3662 = _T_3660_0 & _T_3661_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3664; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3665 = ~_T_3664; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3668; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3669_0; // @[GameUtilities.scala 21:24]
  reg  _T_3669_1; // @[GameUtilities.scala 21:24]
  reg  _T_3670_0; // @[GameUtilities.scala 21:24]
  reg  _T_3670_1; // @[GameUtilities.scala 21:24]
  wire  _T_3671 = _T_3669_0 & _T_3670_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3673; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3674 = ~_T_3673; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3677; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3678_0; // @[GameUtilities.scala 21:24]
  reg  _T_3678_1; // @[GameUtilities.scala 21:24]
  reg  _T_3679_0; // @[GameUtilities.scala 21:24]
  reg  _T_3679_1; // @[GameUtilities.scala 21:24]
  wire  _T_3680 = _T_3678_0 & _T_3679_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3682; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3683 = ~_T_3682; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3686; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3687_0; // @[GameUtilities.scala 21:24]
  reg  _T_3687_1; // @[GameUtilities.scala 21:24]
  reg  _T_3688_0; // @[GameUtilities.scala 21:24]
  reg  _T_3688_1; // @[GameUtilities.scala 21:24]
  wire  _T_3689 = _T_3687_0 & _T_3688_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3691; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3692 = ~_T_3691; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3695; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3696_0; // @[GameUtilities.scala 21:24]
  reg  _T_3696_1; // @[GameUtilities.scala 21:24]
  reg  _T_3697_0; // @[GameUtilities.scala 21:24]
  reg  _T_3697_1; // @[GameUtilities.scala 21:24]
  wire  _T_3698 = _T_3696_0 & _T_3697_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3700; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3701 = ~_T_3700; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3704; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3705_0; // @[GameUtilities.scala 21:24]
  reg  _T_3705_1; // @[GameUtilities.scala 21:24]
  reg  _T_3706_0; // @[GameUtilities.scala 21:24]
  reg  _T_3706_1; // @[GameUtilities.scala 21:24]
  wire  _T_3707 = _T_3705_0 & _T_3706_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3709; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3710 = ~_T_3709; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3713; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3714_0; // @[GameUtilities.scala 21:24]
  reg  _T_3714_1; // @[GameUtilities.scala 21:24]
  reg  _T_3715_0; // @[GameUtilities.scala 21:24]
  reg  _T_3715_1; // @[GameUtilities.scala 21:24]
  wire  _T_3716 = _T_3714_0 & _T_3715_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3718; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3719 = ~_T_3718; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3722; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3723_0; // @[GameUtilities.scala 21:24]
  reg  _T_3723_1; // @[GameUtilities.scala 21:24]
  reg  _T_3724_0; // @[GameUtilities.scala 21:24]
  reg  _T_3724_1; // @[GameUtilities.scala 21:24]
  wire  _T_3725 = _T_3723_0 & _T_3724_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3727; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3728 = ~_T_3727; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3731; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3732_0; // @[GameUtilities.scala 21:24]
  reg  _T_3732_1; // @[GameUtilities.scala 21:24]
  reg  _T_3733_0; // @[GameUtilities.scala 21:24]
  reg  _T_3733_1; // @[GameUtilities.scala 21:24]
  wire  _T_3734 = _T_3732_0 & _T_3733_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3736; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3737 = ~_T_3736; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3740; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3741_0; // @[GameUtilities.scala 21:24]
  reg  _T_3741_1; // @[GameUtilities.scala 21:24]
  reg  _T_3742_0; // @[GameUtilities.scala 21:24]
  reg  _T_3742_1; // @[GameUtilities.scala 21:24]
  wire  _T_3743 = _T_3741_0 & _T_3742_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3745; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3746 = ~_T_3745; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3749; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3750_0; // @[GameUtilities.scala 21:24]
  reg  _T_3750_1; // @[GameUtilities.scala 21:24]
  reg  _T_3751_0; // @[GameUtilities.scala 21:24]
  reg  _T_3751_1; // @[GameUtilities.scala 21:24]
  wire  _T_3752 = _T_3750_0 & _T_3751_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3754; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3755 = ~_T_3754; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3758; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3759_0; // @[GameUtilities.scala 21:24]
  reg  _T_3759_1; // @[GameUtilities.scala 21:24]
  reg  _T_3760_0; // @[GameUtilities.scala 21:24]
  reg  _T_3760_1; // @[GameUtilities.scala 21:24]
  wire  _T_3761 = _T_3759_0 & _T_3760_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3763; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3764 = ~_T_3763; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3767; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3768_0; // @[GameUtilities.scala 21:24]
  reg  _T_3768_1; // @[GameUtilities.scala 21:24]
  reg  _T_3769_0; // @[GameUtilities.scala 21:24]
  reg  _T_3769_1; // @[GameUtilities.scala 21:24]
  wire  _T_3770 = _T_3768_0 & _T_3769_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3772; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3773 = ~_T_3772; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3776; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3777_0; // @[GameUtilities.scala 21:24]
  reg  _T_3777_1; // @[GameUtilities.scala 21:24]
  reg  _T_3778_0; // @[GameUtilities.scala 21:24]
  reg  _T_3778_1; // @[GameUtilities.scala 21:24]
  wire  _T_3779 = _T_3777_0 & _T_3778_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3781; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3782 = ~_T_3781; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3785; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3786_0; // @[GameUtilities.scala 21:24]
  reg  _T_3786_1; // @[GameUtilities.scala 21:24]
  reg  _T_3787_0; // @[GameUtilities.scala 21:24]
  reg  _T_3787_1; // @[GameUtilities.scala 21:24]
  wire  _T_3788 = _T_3786_0 & _T_3787_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3790; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3791 = ~_T_3790; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3794; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3795_0; // @[GameUtilities.scala 21:24]
  reg  _T_3795_1; // @[GameUtilities.scala 21:24]
  reg  _T_3796_0; // @[GameUtilities.scala 21:24]
  reg  _T_3796_1; // @[GameUtilities.scala 21:24]
  wire  _T_3797 = _T_3795_0 & _T_3796_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3799; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3800 = ~_T_3799; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3803; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3805_0; // @[GameUtilities.scala 21:24]
  reg  _T_3805_1; // @[GameUtilities.scala 21:24]
  reg  _T_3808; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3809 = ~_T_3808; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3812; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3814_0; // @[GameUtilities.scala 21:24]
  reg  _T_3814_1; // @[GameUtilities.scala 21:24]
  reg  _T_3817; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3818 = ~_T_3817; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3821; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3823_0; // @[GameUtilities.scala 21:24]
  reg  _T_3823_1; // @[GameUtilities.scala 21:24]
  reg  _T_3826; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3827 = ~_T_3826; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3830; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3832_0; // @[GameUtilities.scala 21:24]
  reg  _T_3832_1; // @[GameUtilities.scala 21:24]
  reg  _T_3835; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3836 = ~_T_3835; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3839; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3841_0; // @[GameUtilities.scala 21:24]
  reg  _T_3841_1; // @[GameUtilities.scala 21:24]
  reg  _T_3844; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3845 = ~_T_3844; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3848; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3850_0; // @[GameUtilities.scala 21:24]
  reg  _T_3850_1; // @[GameUtilities.scala 21:24]
  reg  _T_3853; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3854 = ~_T_3853; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3857; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3859_0; // @[GameUtilities.scala 21:24]
  reg  _T_3859_1; // @[GameUtilities.scala 21:24]
  reg  _T_3862; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3863 = ~_T_3862; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3866; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3867_0; // @[GameUtilities.scala 21:24]
  reg  _T_3867_1; // @[GameUtilities.scala 21:24]
  reg  _T_3868_0; // @[GameUtilities.scala 21:24]
  reg  _T_3868_1; // @[GameUtilities.scala 21:24]
  wire  _T_3869 = _T_3867_0 & _T_3868_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3871; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3872 = ~_T_3871; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3875; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3876_0; // @[GameUtilities.scala 21:24]
  reg  _T_3876_1; // @[GameUtilities.scala 21:24]
  reg  _T_3877_0; // @[GameUtilities.scala 21:24]
  reg  _T_3877_1; // @[GameUtilities.scala 21:24]
  wire  _T_3878 = _T_3876_0 & _T_3877_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3880; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3881 = ~_T_3880; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3884; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3885_0; // @[GameUtilities.scala 21:24]
  reg  _T_3885_1; // @[GameUtilities.scala 21:24]
  reg  _T_3886_0; // @[GameUtilities.scala 21:24]
  reg  _T_3886_1; // @[GameUtilities.scala 21:24]
  wire  _T_3887 = _T_3885_0 & _T_3886_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3889; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3890 = ~_T_3889; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3893; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3894_0; // @[GameUtilities.scala 21:24]
  reg  _T_3894_1; // @[GameUtilities.scala 21:24]
  reg  _T_3895_0; // @[GameUtilities.scala 21:24]
  reg  _T_3895_1; // @[GameUtilities.scala 21:24]
  wire  _T_3896 = _T_3894_0 & _T_3895_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3898; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3899 = ~_T_3898; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3902; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3903_0; // @[GameUtilities.scala 21:24]
  reg  _T_3903_1; // @[GameUtilities.scala 21:24]
  reg  _T_3904_0; // @[GameUtilities.scala 21:24]
  reg  _T_3904_1; // @[GameUtilities.scala 21:24]
  wire  _T_3905 = _T_3903_0 & _T_3904_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3907; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3908 = ~_T_3907; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3911; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3912_0; // @[GameUtilities.scala 21:24]
  reg  _T_3912_1; // @[GameUtilities.scala 21:24]
  reg  _T_3913_0; // @[GameUtilities.scala 21:24]
  reg  _T_3913_1; // @[GameUtilities.scala 21:24]
  wire  _T_3914 = _T_3912_0 & _T_3913_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3916; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3917 = ~_T_3916; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3920; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3921_0; // @[GameUtilities.scala 21:24]
  reg  _T_3921_1; // @[GameUtilities.scala 21:24]
  reg  _T_3922_0; // @[GameUtilities.scala 21:24]
  reg  _T_3922_1; // @[GameUtilities.scala 21:24]
  wire  _T_3923 = _T_3921_0 & _T_3922_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3925; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3926 = ~_T_3925; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3929; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3930_0; // @[GameUtilities.scala 21:24]
  reg  _T_3930_1; // @[GameUtilities.scala 21:24]
  reg  _T_3931_0; // @[GameUtilities.scala 21:24]
  reg  _T_3931_1; // @[GameUtilities.scala 21:24]
  wire  _T_3932 = _T_3930_0 & _T_3931_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3934; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3935 = ~_T_3934; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3938; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3939_0; // @[GameUtilities.scala 21:24]
  reg  _T_3939_1; // @[GameUtilities.scala 21:24]
  reg  _T_3940_0; // @[GameUtilities.scala 21:24]
  reg  _T_3940_1; // @[GameUtilities.scala 21:24]
  wire  _T_3941 = _T_3939_0 & _T_3940_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3943; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3944 = ~_T_3943; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3947; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3948_0; // @[GameUtilities.scala 21:24]
  reg  _T_3948_1; // @[GameUtilities.scala 21:24]
  reg  _T_3949_0; // @[GameUtilities.scala 21:24]
  reg  _T_3949_1; // @[GameUtilities.scala 21:24]
  wire  _T_3950 = _T_3948_0 & _T_3949_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3952; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3953 = ~_T_3952; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3956; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3957_0; // @[GameUtilities.scala 21:24]
  reg  _T_3957_1; // @[GameUtilities.scala 21:24]
  reg  _T_3958_0; // @[GameUtilities.scala 21:24]
  reg  _T_3958_1; // @[GameUtilities.scala 21:24]
  wire  _T_3959 = _T_3957_0 & _T_3958_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3961; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3962 = ~_T_3961; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3965; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3967_0; // @[GameUtilities.scala 21:24]
  reg  _T_3967_1; // @[GameUtilities.scala 21:24]
  reg  _T_3970; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3971 = ~_T_3970; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3974; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3976_0; // @[GameUtilities.scala 21:24]
  reg  _T_3976_1; // @[GameUtilities.scala 21:24]
  reg  _T_3979; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3980 = ~_T_3979; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3983; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3985_0; // @[GameUtilities.scala 21:24]
  reg  _T_3985_1; // @[GameUtilities.scala 21:24]
  reg  _T_3988; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3989 = ~_T_3988; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_3992; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_3993_0; // @[GameUtilities.scala 21:24]
  reg  _T_3993_1; // @[GameUtilities.scala 21:24]
  reg  _T_3994_0; // @[GameUtilities.scala 21:24]
  reg  _T_3994_1; // @[GameUtilities.scala 21:24]
  wire  _T_3995 = _T_3993_0 & _T_3994_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_3997; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_3998 = ~_T_3997; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4001; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4002_0; // @[GameUtilities.scala 21:24]
  reg  _T_4002_1; // @[GameUtilities.scala 21:24]
  reg  _T_4003_0; // @[GameUtilities.scala 21:24]
  reg  _T_4003_1; // @[GameUtilities.scala 21:24]
  wire  _T_4004 = _T_4002_0 & _T_4003_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4006; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4007 = ~_T_4006; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4010; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4011_0; // @[GameUtilities.scala 21:24]
  reg  _T_4011_1; // @[GameUtilities.scala 21:24]
  reg  _T_4012_0; // @[GameUtilities.scala 21:24]
  reg  _T_4012_1; // @[GameUtilities.scala 21:24]
  wire  _T_4013 = _T_4011_0 & _T_4012_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4015; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4016 = ~_T_4015; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4019; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4021_0; // @[GameUtilities.scala 21:24]
  reg  _T_4021_1; // @[GameUtilities.scala 21:24]
  reg  _T_4024; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4025 = ~_T_4024; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4028; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4030_0; // @[GameUtilities.scala 21:24]
  reg  _T_4030_1; // @[GameUtilities.scala 21:24]
  reg  _T_4033; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4034 = ~_T_4033; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4037; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4039_0; // @[GameUtilities.scala 21:24]
  reg  _T_4039_1; // @[GameUtilities.scala 21:24]
  reg  _T_4042; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4043 = ~_T_4042; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4046; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4047_0; // @[GameUtilities.scala 21:24]
  reg  _T_4047_1; // @[GameUtilities.scala 21:24]
  reg  _T_4048_0; // @[GameUtilities.scala 21:24]
  reg  _T_4048_1; // @[GameUtilities.scala 21:24]
  wire  _T_4049 = _T_4047_0 & _T_4048_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4051; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4052 = ~_T_4051; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4055; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4056_0; // @[GameUtilities.scala 21:24]
  reg  _T_4056_1; // @[GameUtilities.scala 21:24]
  reg  _T_4057_0; // @[GameUtilities.scala 21:24]
  reg  _T_4057_1; // @[GameUtilities.scala 21:24]
  wire  _T_4058 = _T_4056_0 & _T_4057_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4060; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4061 = ~_T_4060; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4064; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4065_0; // @[GameUtilities.scala 21:24]
  reg  _T_4065_1; // @[GameUtilities.scala 21:24]
  reg  _T_4066_0; // @[GameUtilities.scala 21:24]
  reg  _T_4066_1; // @[GameUtilities.scala 21:24]
  wire  _T_4067 = _T_4065_0 & _T_4066_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4069; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4070 = ~_T_4069; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4073; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4074_0; // @[GameUtilities.scala 21:24]
  reg  _T_4074_1; // @[GameUtilities.scala 21:24]
  reg  _T_4075_0; // @[GameUtilities.scala 21:24]
  reg  _T_4075_1; // @[GameUtilities.scala 21:24]
  wire  _T_4076 = _T_4074_0 & _T_4075_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4078; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4079 = ~_T_4078; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4082; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4083_0; // @[GameUtilities.scala 21:24]
  reg  _T_4083_1; // @[GameUtilities.scala 21:24]
  reg  _T_4084_0; // @[GameUtilities.scala 21:24]
  reg  _T_4084_1; // @[GameUtilities.scala 21:24]
  wire  _T_4085 = _T_4083_0 & _T_4084_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4087; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4088 = ~_T_4087; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4091; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4092_0; // @[GameUtilities.scala 21:24]
  reg  _T_4092_1; // @[GameUtilities.scala 21:24]
  reg  _T_4093_0; // @[GameUtilities.scala 21:24]
  reg  _T_4093_1; // @[GameUtilities.scala 21:24]
  wire  _T_4094 = _T_4092_0 & _T_4093_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4096; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4097 = ~_T_4096; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4100; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4102_0; // @[GameUtilities.scala 21:24]
  reg  _T_4102_1; // @[GameUtilities.scala 21:24]
  reg  _T_4105; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4106 = ~_T_4105; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4109; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4111_0; // @[GameUtilities.scala 21:24]
  reg  _T_4111_1; // @[GameUtilities.scala 21:24]
  reg  _T_4114; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4115 = ~_T_4114; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4118; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4120_0; // @[GameUtilities.scala 21:24]
  reg  _T_4120_1; // @[GameUtilities.scala 21:24]
  reg  _T_4123; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4124 = ~_T_4123; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4127; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4128_0; // @[GameUtilities.scala 21:24]
  reg  _T_4128_1; // @[GameUtilities.scala 21:24]
  reg  _T_4129_0; // @[GameUtilities.scala 21:24]
  reg  _T_4129_1; // @[GameUtilities.scala 21:24]
  wire  _T_4130 = _T_4128_0 & _T_4129_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4132; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4133 = ~_T_4132; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4136; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4137_0; // @[GameUtilities.scala 21:24]
  reg  _T_4137_1; // @[GameUtilities.scala 21:24]
  reg  _T_4138_0; // @[GameUtilities.scala 21:24]
  reg  _T_4138_1; // @[GameUtilities.scala 21:24]
  wire  _T_4139 = _T_4137_0 & _T_4138_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4141; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4142 = ~_T_4141; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4145; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4146_0; // @[GameUtilities.scala 21:24]
  reg  _T_4146_1; // @[GameUtilities.scala 21:24]
  reg  _T_4147_0; // @[GameUtilities.scala 21:24]
  reg  _T_4147_1; // @[GameUtilities.scala 21:24]
  wire  _T_4148 = _T_4146_0 & _T_4147_0; // @[GraphicEngineVGA.scala 309:91]
  reg  _T_4150; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4151 = ~_T_4150; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4154; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4156_0; // @[GameUtilities.scala 21:24]
  reg  _T_4156_1; // @[GameUtilities.scala 21:24]
  reg  _T_4159; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4160 = ~_T_4159; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4163; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4165_0; // @[GameUtilities.scala 21:24]
  reg  _T_4165_1; // @[GameUtilities.scala 21:24]
  reg  _T_4168; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4169 = ~_T_4168; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4172; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4174_0; // @[GameUtilities.scala 21:24]
  reg  _T_4174_1; // @[GameUtilities.scala 21:24]
  reg  _T_4177; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4178 = ~_T_4177; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4181; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4183_0; // @[GameUtilities.scala 21:24]
  reg  _T_4183_1; // @[GameUtilities.scala 21:24]
  reg  _T_4186; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4187 = ~_T_4186; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4190; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4192_0; // @[GameUtilities.scala 21:24]
  reg  _T_4192_1; // @[GameUtilities.scala 21:24]
  reg  _T_4195; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4196 = ~_T_4195; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4199; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4201_0; // @[GameUtilities.scala 21:24]
  reg  _T_4201_1; // @[GameUtilities.scala 21:24]
  reg  _T_4204; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4205 = ~_T_4204; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4208; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4210_0; // @[GameUtilities.scala 21:24]
  reg  _T_4210_1; // @[GameUtilities.scala 21:24]
  reg  _T_4213; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4214 = ~_T_4213; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4217; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4219_0; // @[GameUtilities.scala 21:24]
  reg  _T_4219_1; // @[GameUtilities.scala 21:24]
  reg  _T_4222; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4223 = ~_T_4222; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4226; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4228_0; // @[GameUtilities.scala 21:24]
  reg  _T_4228_1; // @[GameUtilities.scala 21:24]
  reg  _T_4231; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4232 = ~_T_4231; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4235; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4237_0; // @[GameUtilities.scala 21:24]
  reg  _T_4237_1; // @[GameUtilities.scala 21:24]
  reg  _T_4240; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4241 = ~_T_4240; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4244; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4246_0; // @[GameUtilities.scala 21:24]
  reg  _T_4246_1; // @[GameUtilities.scala 21:24]
  reg  _T_4249; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4250 = ~_T_4249; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4253; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4255_0; // @[GameUtilities.scala 21:24]
  reg  _T_4255_1; // @[GameUtilities.scala 21:24]
  reg  _T_4258; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4259 = ~_T_4258; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4262; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4264_0; // @[GameUtilities.scala 21:24]
  reg  _T_4264_1; // @[GameUtilities.scala 21:24]
  reg  _T_4267; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4268 = ~_T_4267; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4271; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4273_0; // @[GameUtilities.scala 21:24]
  reg  _T_4273_1; // @[GameUtilities.scala 21:24]
  reg  _T_4276; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4277 = ~_T_4276; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4280; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4282_0; // @[GameUtilities.scala 21:24]
  reg  _T_4282_1; // @[GameUtilities.scala 21:24]
  reg  _T_4285; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4286 = ~_T_4285; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4289; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4291_0; // @[GameUtilities.scala 21:24]
  reg  _T_4291_1; // @[GameUtilities.scala 21:24]
  reg  _T_4294; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4295 = ~_T_4294; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4298; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4300_0; // @[GameUtilities.scala 21:24]
  reg  _T_4300_1; // @[GameUtilities.scala 21:24]
  reg  _T_4303; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4304 = ~_T_4303; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4307; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4309_0; // @[GameUtilities.scala 21:24]
  reg  _T_4309_1; // @[GameUtilities.scala 21:24]
  reg  _T_4312; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4313 = ~_T_4312; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4316; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4318_0; // @[GameUtilities.scala 21:24]
  reg  _T_4318_1; // @[GameUtilities.scala 21:24]
  reg  _T_4321; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4322 = ~_T_4321; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4325; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4327_0; // @[GameUtilities.scala 21:24]
  reg  _T_4327_1; // @[GameUtilities.scala 21:24]
  reg  _T_4330; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4331 = ~_T_4330; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4334; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4336_0; // @[GameUtilities.scala 21:24]
  reg  _T_4336_1; // @[GameUtilities.scala 21:24]
  reg  _T_4339; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4340 = ~_T_4339; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4343; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4345_0; // @[GameUtilities.scala 21:24]
  reg  _T_4345_1; // @[GameUtilities.scala 21:24]
  reg  _T_4348; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4349 = ~_T_4348; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4352; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4354_0; // @[GameUtilities.scala 21:24]
  reg  _T_4354_1; // @[GameUtilities.scala 21:24]
  reg  _T_4357; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4358 = ~_T_4357; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4361; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4363_0; // @[GameUtilities.scala 21:24]
  reg  _T_4363_1; // @[GameUtilities.scala 21:24]
  reg  _T_4366; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4367 = ~_T_4366; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4370; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4372_0; // @[GameUtilities.scala 21:24]
  reg  _T_4372_1; // @[GameUtilities.scala 21:24]
  reg  _T_4375; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4376 = ~_T_4375; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4379; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4381_0; // @[GameUtilities.scala 21:24]
  reg  _T_4381_1; // @[GameUtilities.scala 21:24]
  reg  _T_4384; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4385 = ~_T_4384; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4388; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4390_0; // @[GameUtilities.scala 21:24]
  reg  _T_4390_1; // @[GameUtilities.scala 21:24]
  reg  _T_4393; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4394 = ~_T_4393; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4397; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4399_0; // @[GameUtilities.scala 21:24]
  reg  _T_4399_1; // @[GameUtilities.scala 21:24]
  reg  _T_4402; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4403 = ~_T_4402; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4406; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4408_0; // @[GameUtilities.scala 21:24]
  reg  _T_4408_1; // @[GameUtilities.scala 21:24]
  reg  _T_4411; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4412 = ~_T_4411; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4415; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4417_0; // @[GameUtilities.scala 21:24]
  reg  _T_4417_1; // @[GameUtilities.scala 21:24]
  reg  _T_4420; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4421 = ~_T_4420; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4424; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4426_0; // @[GameUtilities.scala 21:24]
  reg  _T_4426_1; // @[GameUtilities.scala 21:24]
  reg  _T_4429; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4430 = ~_T_4429; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4433; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4435_0; // @[GameUtilities.scala 21:24]
  reg  _T_4435_1; // @[GameUtilities.scala 21:24]
  reg  _T_4438; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4439 = ~_T_4438; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4442; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4444_0; // @[GameUtilities.scala 21:24]
  reg  _T_4444_1; // @[GameUtilities.scala 21:24]
  reg  _T_4447; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4448 = ~_T_4447; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4451; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4453_0; // @[GameUtilities.scala 21:24]
  reg  _T_4453_1; // @[GameUtilities.scala 21:24]
  reg  _T_4456; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4457 = ~_T_4456; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4460; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4462_0; // @[GameUtilities.scala 21:24]
  reg  _T_4462_1; // @[GameUtilities.scala 21:24]
  reg  _T_4465; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4466 = ~_T_4465; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4469; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4471_0; // @[GameUtilities.scala 21:24]
  reg  _T_4471_1; // @[GameUtilities.scala 21:24]
  reg  _T_4474; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4475 = ~_T_4474; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4478; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4480_0; // @[GameUtilities.scala 21:24]
  reg  _T_4480_1; // @[GameUtilities.scala 21:24]
  reg  _T_4483; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4484 = ~_T_4483; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4487; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4489_0; // @[GameUtilities.scala 21:24]
  reg  _T_4489_1; // @[GameUtilities.scala 21:24]
  reg  _T_4492; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4493 = ~_T_4492; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4496; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4498_0; // @[GameUtilities.scala 21:24]
  reg  _T_4498_1; // @[GameUtilities.scala 21:24]
  reg  _T_4501; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4502 = ~_T_4501; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4505; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4507_0; // @[GameUtilities.scala 21:24]
  reg  _T_4507_1; // @[GameUtilities.scala 21:24]
  reg  _T_4510; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4511 = ~_T_4510; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4514; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4516_0; // @[GameUtilities.scala 21:24]
  reg  _T_4516_1; // @[GameUtilities.scala 21:24]
  reg  _T_4519; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4520 = ~_T_4519; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4523; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4525_0; // @[GameUtilities.scala 21:24]
  reg  _T_4525_1; // @[GameUtilities.scala 21:24]
  reg  _T_4528; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4529 = ~_T_4528; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4532; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4534_0; // @[GameUtilities.scala 21:24]
  reg  _T_4534_1; // @[GameUtilities.scala 21:24]
  reg  _T_4537; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4538 = ~_T_4537; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4541; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4543_0; // @[GameUtilities.scala 21:24]
  reg  _T_4543_1; // @[GameUtilities.scala 21:24]
  reg  _T_4546; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4547 = ~_T_4546; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4550; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4552_0; // @[GameUtilities.scala 21:24]
  reg  _T_4552_1; // @[GameUtilities.scala 21:24]
  reg  _T_4555; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4556 = ~_T_4555; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4559; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4561_0; // @[GameUtilities.scala 21:24]
  reg  _T_4561_1; // @[GameUtilities.scala 21:24]
  reg  _T_4564; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4565 = ~_T_4564; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4568; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4570_0; // @[GameUtilities.scala 21:24]
  reg  _T_4570_1; // @[GameUtilities.scala 21:24]
  reg  _T_4573; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4574 = ~_T_4573; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4577; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4579_0; // @[GameUtilities.scala 21:24]
  reg  _T_4579_1; // @[GameUtilities.scala 21:24]
  reg  _T_4582; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4583 = ~_T_4582; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4586; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4588_0; // @[GameUtilities.scala 21:24]
  reg  _T_4588_1; // @[GameUtilities.scala 21:24]
  reg  _T_4591; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4592 = ~_T_4591; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4595; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4597_0; // @[GameUtilities.scala 21:24]
  reg  _T_4597_1; // @[GameUtilities.scala 21:24]
  reg  _T_4600; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4601 = ~_T_4600; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4604; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4606_0; // @[GameUtilities.scala 21:24]
  reg  _T_4606_1; // @[GameUtilities.scala 21:24]
  reg  _T_4609; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4610 = ~_T_4609; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4613; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4615_0; // @[GameUtilities.scala 21:24]
  reg  _T_4615_1; // @[GameUtilities.scala 21:24]
  reg  _T_4618; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4619 = ~_T_4618; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4622; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4624_0; // @[GameUtilities.scala 21:24]
  reg  _T_4624_1; // @[GameUtilities.scala 21:24]
  reg  _T_4627; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4628 = ~_T_4627; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4631; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4633_0; // @[GameUtilities.scala 21:24]
  reg  _T_4633_1; // @[GameUtilities.scala 21:24]
  reg  _T_4636; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4637 = ~_T_4636; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] _T_4640; // @[GraphicEngineVGA.scala 308:60]
  reg  _T_4642_0; // @[GameUtilities.scala 21:24]
  reg  _T_4642_1; // @[GameUtilities.scala 21:24]
  reg  _T_4645; // @[GraphicEngineVGA.scala 309:132]
  wire  _T_4646 = ~_T_4645; // @[GraphicEngineVGA.scala 309:123]
  reg [5:0] pixelColorSprite; // @[GraphicEngineVGA.scala 311:33]
  reg  pixelColorSpriteValid; // @[GraphicEngineVGA.scala 312:38]
  wire [5:0] pixelColorInDisplay = pixelColorSpriteValid ? pixelColorSprite : pixelColorBack; // @[GraphicEngineVGA.scala 316:32]
  reg  _T_4648_0; // @[GameUtilities.scala 21:24]
  reg  _T_4648_1; // @[GameUtilities.scala 21:24]
  reg  _T_4648_2; // @[GameUtilities.scala 21:24]
  wire [5:0] pixelColourVGA = _T_4648_0 ? pixelColorInDisplay : 6'h0; // @[GraphicEngineVGA.scala 317:27]
  reg [3:0] _T_4655; // @[GraphicEngineVGA.scala 321:23]
  reg [3:0] _T_4656; // @[GraphicEngineVGA.scala 322:25]
  reg [3:0] _T_4657; // @[GraphicEngineVGA.scala 323:24]
  Memory backTileMemories_0_0 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_0_clock),
    .io_address(backTileMemories_0_0_io_address),
    .io_dataRead(backTileMemories_0_0_io_dataRead)
  );
  Memory_1 backTileMemories_0_1 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_1_clock),
    .io_address(backTileMemories_0_1_io_address),
    .io_dataRead(backTileMemories_0_1_io_dataRead)
  );
  Memory_2 backTileMemories_0_2 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_2_clock),
    .io_address(backTileMemories_0_2_io_address),
    .io_dataRead(backTileMemories_0_2_io_dataRead)
  );
  Memory_3 backTileMemories_0_3 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_3_clock),
    .io_address(backTileMemories_0_3_io_address),
    .io_dataRead(backTileMemories_0_3_io_dataRead)
  );
  Memory_4 backTileMemories_0_4 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_4_clock),
    .io_address(backTileMemories_0_4_io_address),
    .io_dataRead(backTileMemories_0_4_io_dataRead)
  );
  Memory_5 backTileMemories_0_5 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_5_clock),
    .io_address(backTileMemories_0_5_io_address),
    .io_dataRead(backTileMemories_0_5_io_dataRead)
  );
  Memory_6 backTileMemories_0_6 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_6_clock),
    .io_address(backTileMemories_0_6_io_address),
    .io_dataRead(backTileMemories_0_6_io_dataRead)
  );
  Memory_7 backTileMemories_0_7 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_7_clock),
    .io_address(backTileMemories_0_7_io_address),
    .io_dataRead(backTileMemories_0_7_io_dataRead)
  );
  Memory_8 backTileMemories_0_8 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_8_clock),
    .io_address(backTileMemories_0_8_io_address),
    .io_dataRead(backTileMemories_0_8_io_dataRead)
  );
  Memory_9 backTileMemories_0_9 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_9_clock),
    .io_address(backTileMemories_0_9_io_address),
    .io_dataRead(backTileMemories_0_9_io_dataRead)
  );
  Memory_10 backTileMemories_0_10 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_10_clock),
    .io_address(backTileMemories_0_10_io_address),
    .io_dataRead(backTileMemories_0_10_io_dataRead)
  );
  Memory_11 backTileMemories_0_11 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_11_clock),
    .io_address(backTileMemories_0_11_io_address),
    .io_dataRead(backTileMemories_0_11_io_dataRead)
  );
  Memory_12 backTileMemories_0_12 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_12_clock),
    .io_address(backTileMemories_0_12_io_address),
    .io_dataRead(backTileMemories_0_12_io_dataRead)
  );
  Memory_13 backTileMemories_0_13 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_13_clock),
    .io_address(backTileMemories_0_13_io_address),
    .io_dataRead(backTileMemories_0_13_io_dataRead)
  );
  Memory_14 backTileMemories_0_14 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_14_clock),
    .io_address(backTileMemories_0_14_io_address),
    .io_dataRead(backTileMemories_0_14_io_dataRead)
  );
  Memory_15 backTileMemories_0_15 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_15_clock),
    .io_address(backTileMemories_0_15_io_address),
    .io_dataRead(backTileMemories_0_15_io_dataRead)
  );
  Memory_16 backTileMemories_0_16 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_16_clock),
    .io_address(backTileMemories_0_16_io_address),
    .io_dataRead(backTileMemories_0_16_io_dataRead)
  );
  Memory_17 backTileMemories_0_17 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_17_clock),
    .io_address(backTileMemories_0_17_io_address),
    .io_dataRead(backTileMemories_0_17_io_dataRead)
  );
  Memory_18 backTileMemories_0_18 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_18_clock),
    .io_address(backTileMemories_0_18_io_address),
    .io_dataRead(backTileMemories_0_18_io_dataRead)
  );
  Memory_19 backTileMemories_0_19 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_19_clock),
    .io_address(backTileMemories_0_19_io_address),
    .io_dataRead(backTileMemories_0_19_io_dataRead)
  );
  Memory_20 backTileMemories_0_20 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_20_clock),
    .io_address(backTileMemories_0_20_io_address),
    .io_dataRead(backTileMemories_0_20_io_dataRead)
  );
  Memory_21 backTileMemories_0_21 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_21_clock),
    .io_address(backTileMemories_0_21_io_address),
    .io_dataRead(backTileMemories_0_21_io_dataRead)
  );
  Memory_22 backTileMemories_0_22 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_22_clock),
    .io_address(backTileMemories_0_22_io_address),
    .io_dataRead(backTileMemories_0_22_io_dataRead)
  );
  Memory_23 backTileMemories_0_23 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_23_clock),
    .io_address(backTileMemories_0_23_io_address),
    .io_dataRead(backTileMemories_0_23_io_dataRead)
  );
  Memory_24 backTileMemories_0_24 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_24_clock),
    .io_address(backTileMemories_0_24_io_address),
    .io_dataRead(backTileMemories_0_24_io_dataRead)
  );
  Memory_25 backTileMemories_0_25 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_25_clock),
    .io_address(backTileMemories_0_25_io_address),
    .io_dataRead(backTileMemories_0_25_io_dataRead)
  );
  Memory_26 backTileMemories_0_26 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_26_clock),
    .io_address(backTileMemories_0_26_io_address),
    .io_dataRead(backTileMemories_0_26_io_dataRead)
  );
  Memory_27 backTileMemories_0_27 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_27_clock),
    .io_address(backTileMemories_0_27_io_address),
    .io_dataRead(backTileMemories_0_27_io_dataRead)
  );
  Memory_28 backTileMemories_0_28 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_28_clock),
    .io_address(backTileMemories_0_28_io_address),
    .io_dataRead(backTileMemories_0_28_io_dataRead)
  );
  Memory_29 backTileMemories_0_29 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_29_clock),
    .io_address(backTileMemories_0_29_io_address),
    .io_dataRead(backTileMemories_0_29_io_dataRead)
  );
  Memory_30 backTileMemories_0_30 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_30_clock),
    .io_address(backTileMemories_0_30_io_address),
    .io_dataRead(backTileMemories_0_30_io_dataRead)
  );
  Memory_31 backTileMemories_0_31 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_0_31_clock),
    .io_address(backTileMemories_0_31_io_address),
    .io_dataRead(backTileMemories_0_31_io_dataRead)
  );
  Memory backTileMemories_1_0 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_0_clock),
    .io_address(backTileMemories_1_0_io_address),
    .io_dataRead(backTileMemories_1_0_io_dataRead)
  );
  Memory_1 backTileMemories_1_1 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_1_clock),
    .io_address(backTileMemories_1_1_io_address),
    .io_dataRead(backTileMemories_1_1_io_dataRead)
  );
  Memory_2 backTileMemories_1_2 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_2_clock),
    .io_address(backTileMemories_1_2_io_address),
    .io_dataRead(backTileMemories_1_2_io_dataRead)
  );
  Memory_3 backTileMemories_1_3 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_3_clock),
    .io_address(backTileMemories_1_3_io_address),
    .io_dataRead(backTileMemories_1_3_io_dataRead)
  );
  Memory_4 backTileMemories_1_4 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_4_clock),
    .io_address(backTileMemories_1_4_io_address),
    .io_dataRead(backTileMemories_1_4_io_dataRead)
  );
  Memory_5 backTileMemories_1_5 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_5_clock),
    .io_address(backTileMemories_1_5_io_address),
    .io_dataRead(backTileMemories_1_5_io_dataRead)
  );
  Memory_6 backTileMemories_1_6 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_6_clock),
    .io_address(backTileMemories_1_6_io_address),
    .io_dataRead(backTileMemories_1_6_io_dataRead)
  );
  Memory_7 backTileMemories_1_7 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_7_clock),
    .io_address(backTileMemories_1_7_io_address),
    .io_dataRead(backTileMemories_1_7_io_dataRead)
  );
  Memory_8 backTileMemories_1_8 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_8_clock),
    .io_address(backTileMemories_1_8_io_address),
    .io_dataRead(backTileMemories_1_8_io_dataRead)
  );
  Memory_9 backTileMemories_1_9 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_9_clock),
    .io_address(backTileMemories_1_9_io_address),
    .io_dataRead(backTileMemories_1_9_io_dataRead)
  );
  Memory_10 backTileMemories_1_10 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_10_clock),
    .io_address(backTileMemories_1_10_io_address),
    .io_dataRead(backTileMemories_1_10_io_dataRead)
  );
  Memory_11 backTileMemories_1_11 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_11_clock),
    .io_address(backTileMemories_1_11_io_address),
    .io_dataRead(backTileMemories_1_11_io_dataRead)
  );
  Memory_12 backTileMemories_1_12 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_12_clock),
    .io_address(backTileMemories_1_12_io_address),
    .io_dataRead(backTileMemories_1_12_io_dataRead)
  );
  Memory_13 backTileMemories_1_13 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_13_clock),
    .io_address(backTileMemories_1_13_io_address),
    .io_dataRead(backTileMemories_1_13_io_dataRead)
  );
  Memory_14 backTileMemories_1_14 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_14_clock),
    .io_address(backTileMemories_1_14_io_address),
    .io_dataRead(backTileMemories_1_14_io_dataRead)
  );
  Memory_15 backTileMemories_1_15 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_15_clock),
    .io_address(backTileMemories_1_15_io_address),
    .io_dataRead(backTileMemories_1_15_io_dataRead)
  );
  Memory_16 backTileMemories_1_16 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_16_clock),
    .io_address(backTileMemories_1_16_io_address),
    .io_dataRead(backTileMemories_1_16_io_dataRead)
  );
  Memory_17 backTileMemories_1_17 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_17_clock),
    .io_address(backTileMemories_1_17_io_address),
    .io_dataRead(backTileMemories_1_17_io_dataRead)
  );
  Memory_18 backTileMemories_1_18 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_18_clock),
    .io_address(backTileMemories_1_18_io_address),
    .io_dataRead(backTileMemories_1_18_io_dataRead)
  );
  Memory_19 backTileMemories_1_19 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_19_clock),
    .io_address(backTileMemories_1_19_io_address),
    .io_dataRead(backTileMemories_1_19_io_dataRead)
  );
  Memory_20 backTileMemories_1_20 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_20_clock),
    .io_address(backTileMemories_1_20_io_address),
    .io_dataRead(backTileMemories_1_20_io_dataRead)
  );
  Memory_21 backTileMemories_1_21 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_21_clock),
    .io_address(backTileMemories_1_21_io_address),
    .io_dataRead(backTileMemories_1_21_io_dataRead)
  );
  Memory_22 backTileMemories_1_22 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_22_clock),
    .io_address(backTileMemories_1_22_io_address),
    .io_dataRead(backTileMemories_1_22_io_dataRead)
  );
  Memory_23 backTileMemories_1_23 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_23_clock),
    .io_address(backTileMemories_1_23_io_address),
    .io_dataRead(backTileMemories_1_23_io_dataRead)
  );
  Memory_24 backTileMemories_1_24 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_24_clock),
    .io_address(backTileMemories_1_24_io_address),
    .io_dataRead(backTileMemories_1_24_io_dataRead)
  );
  Memory_25 backTileMemories_1_25 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_25_clock),
    .io_address(backTileMemories_1_25_io_address),
    .io_dataRead(backTileMemories_1_25_io_dataRead)
  );
  Memory_26 backTileMemories_1_26 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_26_clock),
    .io_address(backTileMemories_1_26_io_address),
    .io_dataRead(backTileMemories_1_26_io_dataRead)
  );
  Memory_27 backTileMemories_1_27 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_27_clock),
    .io_address(backTileMemories_1_27_io_address),
    .io_dataRead(backTileMemories_1_27_io_dataRead)
  );
  Memory_28 backTileMemories_1_28 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_28_clock),
    .io_address(backTileMemories_1_28_io_address),
    .io_dataRead(backTileMemories_1_28_io_dataRead)
  );
  Memory_29 backTileMemories_1_29 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_29_clock),
    .io_address(backTileMemories_1_29_io_address),
    .io_dataRead(backTileMemories_1_29_io_dataRead)
  );
  Memory_30 backTileMemories_1_30 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_30_clock),
    .io_address(backTileMemories_1_30_io_address),
    .io_dataRead(backTileMemories_1_30_io_dataRead)
  );
  Memory_31 backTileMemories_1_31 ( // @[GraphicEngineVGA.scala 162:34]
    .clock(backTileMemories_1_31_clock),
    .io_address(backTileMemories_1_31_io_address),
    .io_dataRead(backTileMemories_1_31_io_dataRead)
  );
  Memory_64 backBufferMemories_0 ( // @[GraphicEngineVGA.scala 186:34]
    .clock(backBufferMemories_0_clock),
    .io_address(backBufferMemories_0_io_address),
    .io_dataRead(backBufferMemories_0_io_dataRead),
    .io_writeEnable(backBufferMemories_0_io_writeEnable),
    .io_dataWrite(backBufferMemories_0_io_dataWrite)
  );
  Memory_64 backBufferMemories_1 ( // @[GraphicEngineVGA.scala 186:34]
    .clock(backBufferMemories_1_clock),
    .io_address(backBufferMemories_1_io_address),
    .io_dataRead(backBufferMemories_1_io_dataRead),
    .io_writeEnable(backBufferMemories_1_io_writeEnable),
    .io_dataWrite(backBufferMemories_1_io_dataWrite)
  );
  Memory_64 backBufferShadowMemories_0 ( // @[GraphicEngineVGA.scala 191:40]
    .clock(backBufferShadowMemories_0_clock),
    .io_address(backBufferShadowMemories_0_io_address),
    .io_dataRead(backBufferShadowMemories_0_io_dataRead),
    .io_writeEnable(backBufferShadowMemories_0_io_writeEnable),
    .io_dataWrite(backBufferShadowMemories_0_io_dataWrite)
  );
  Memory_64 backBufferShadowMemories_1 ( // @[GraphicEngineVGA.scala 191:40]
    .clock(backBufferShadowMemories_1_clock),
    .io_address(backBufferShadowMemories_1_io_address),
    .io_dataRead(backBufferShadowMemories_1_io_dataRead),
    .io_writeEnable(backBufferShadowMemories_1_io_writeEnable),
    .io_dataWrite(backBufferShadowMemories_1_io_dataWrite)
  );
  Memory_68 backBufferRestoreMemories_0 ( // @[GraphicEngineVGA.scala 197:41]
    .clock(backBufferRestoreMemories_0_clock),
    .io_address(backBufferRestoreMemories_0_io_address),
    .io_dataRead(backBufferRestoreMemories_0_io_dataRead)
  );
  Memory_69 backBufferRestoreMemories_1 ( // @[GraphicEngineVGA.scala 197:41]
    .clock(backBufferRestoreMemories_1_clock),
    .io_address(backBufferRestoreMemories_1_io_address),
    .io_dataRead(backBufferRestoreMemories_1_io_dataRead)
  );
  Memory_70 spriteMemories_0 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_0_clock),
    .io_address(spriteMemories_0_io_address),
    .io_dataRead(spriteMemories_0_io_dataRead)
  );
  Memory_71 spriteMemories_1 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_1_clock),
    .io_address(spriteMemories_1_io_address),
    .io_dataRead(spriteMemories_1_io_dataRead)
  );
  Memory_72 spriteMemories_2 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_2_clock),
    .io_address(spriteMemories_2_io_address),
    .io_dataRead(spriteMemories_2_io_dataRead)
  );
  Memory_73 spriteMemories_3 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_3_clock),
    .io_address(spriteMemories_3_io_address),
    .io_dataRead(spriteMemories_3_io_dataRead)
  );
  Memory_74 spriteMemories_4 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_4_clock),
    .io_address(spriteMemories_4_io_address),
    .io_dataRead(spriteMemories_4_io_dataRead)
  );
  Memory_75 spriteMemories_5 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_5_clock),
    .io_address(spriteMemories_5_io_address),
    .io_dataRead(spriteMemories_5_io_dataRead)
  );
  Memory_76 spriteMemories_6 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_6_clock),
    .io_address(spriteMemories_6_io_address),
    .io_dataRead(spriteMemories_6_io_dataRead)
  );
  Memory_77 spriteMemories_7 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_7_clock),
    .io_address(spriteMemories_7_io_address),
    .io_dataRead(spriteMemories_7_io_dataRead)
  );
  Memory_78 spriteMemories_8 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_8_clock),
    .io_address(spriteMemories_8_io_address),
    .io_dataRead(spriteMemories_8_io_dataRead)
  );
  Memory_79 spriteMemories_9 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_9_clock),
    .io_address(spriteMemories_9_io_address),
    .io_dataRead(spriteMemories_9_io_dataRead)
  );
  Memory_80 spriteMemories_10 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_10_clock),
    .io_address(spriteMemories_10_io_address),
    .io_dataRead(spriteMemories_10_io_dataRead)
  );
  Memory_81 spriteMemories_11 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_11_clock),
    .io_address(spriteMemories_11_io_address),
    .io_dataRead(spriteMemories_11_io_dataRead)
  );
  Memory_82 spriteMemories_12 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_12_clock),
    .io_address(spriteMemories_12_io_address),
    .io_dataRead(spriteMemories_12_io_dataRead)
  );
  Memory_83 spriteMemories_13 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_13_clock),
    .io_address(spriteMemories_13_io_address),
    .io_dataRead(spriteMemories_13_io_dataRead)
  );
  Memory_84 spriteMemories_14 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_14_clock),
    .io_address(spriteMemories_14_io_address),
    .io_dataRead(spriteMemories_14_io_dataRead)
  );
  Memory_85 spriteMemories_15 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_15_clock),
    .io_address(spriteMemories_15_io_address),
    .io_dataRead(spriteMemories_15_io_dataRead)
  );
  Memory_86 spriteMemories_16 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_16_clock),
    .io_address(spriteMemories_16_io_address),
    .io_dataRead(spriteMemories_16_io_dataRead)
  );
  Memory_87 spriteMemories_17 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_17_clock),
    .io_address(spriteMemories_17_io_address),
    .io_dataRead(spriteMemories_17_io_dataRead)
  );
  Memory_88 spriteMemories_18 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_18_clock),
    .io_address(spriteMemories_18_io_address),
    .io_dataRead(spriteMemories_18_io_dataRead)
  );
  Memory_89 spriteMemories_19 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_19_clock),
    .io_address(spriteMemories_19_io_address),
    .io_dataRead(spriteMemories_19_io_dataRead)
  );
  Memory_90 spriteMemories_20 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_20_clock),
    .io_address(spriteMemories_20_io_address),
    .io_dataRead(spriteMemories_20_io_dataRead)
  );
  Memory_91 spriteMemories_21 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_21_clock),
    .io_address(spriteMemories_21_io_address),
    .io_dataRead(spriteMemories_21_io_dataRead)
  );
  Memory_92 spriteMemories_22 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_22_clock),
    .io_address(spriteMemories_22_io_address),
    .io_dataRead(spriteMemories_22_io_dataRead)
  );
  Memory_93 spriteMemories_23 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_23_clock),
    .io_address(spriteMemories_23_io_address),
    .io_dataRead(spriteMemories_23_io_dataRead)
  );
  Memory_94 spriteMemories_24 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_24_clock),
    .io_address(spriteMemories_24_io_address),
    .io_dataRead(spriteMemories_24_io_dataRead)
  );
  Memory_95 spriteMemories_25 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_25_clock),
    .io_address(spriteMemories_25_io_address),
    .io_dataRead(spriteMemories_25_io_dataRead)
  );
  Memory_96 spriteMemories_26 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_26_clock),
    .io_address(spriteMemories_26_io_address),
    .io_dataRead(spriteMemories_26_io_dataRead)
  );
  Memory_97 spriteMemories_27 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_27_clock),
    .io_address(spriteMemories_27_io_address),
    .io_dataRead(spriteMemories_27_io_dataRead)
  );
  Memory_98 spriteMemories_28 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_28_clock),
    .io_address(spriteMemories_28_io_address),
    .io_dataRead(spriteMemories_28_io_dataRead)
  );
  Memory_99 spriteMemories_29 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_29_clock),
    .io_address(spriteMemories_29_io_address),
    .io_dataRead(spriteMemories_29_io_dataRead)
  );
  Memory_100 spriteMemories_30 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_30_clock),
    .io_address(spriteMemories_30_io_address),
    .io_dataRead(spriteMemories_30_io_dataRead)
  );
  Memory_101 spriteMemories_31 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_31_clock),
    .io_address(spriteMemories_31_io_address),
    .io_dataRead(spriteMemories_31_io_dataRead)
  );
  Memory_102 spriteMemories_32 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_32_clock),
    .io_address(spriteMemories_32_io_address),
    .io_dataRead(spriteMemories_32_io_dataRead)
  );
  Memory_103 spriteMemories_33 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_33_clock),
    .io_address(spriteMemories_33_io_address),
    .io_dataRead(spriteMemories_33_io_dataRead)
  );
  Memory_104 spriteMemories_34 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_34_clock),
    .io_address(spriteMemories_34_io_address),
    .io_dataRead(spriteMemories_34_io_dataRead)
  );
  Memory_105 spriteMemories_35 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_35_clock),
    .io_address(spriteMemories_35_io_address),
    .io_dataRead(spriteMemories_35_io_dataRead)
  );
  Memory_106 spriteMemories_36 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_36_clock),
    .io_address(spriteMemories_36_io_address),
    .io_dataRead(spriteMemories_36_io_dataRead)
  );
  Memory_107 spriteMemories_37 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_37_clock),
    .io_address(spriteMemories_37_io_address),
    .io_dataRead(spriteMemories_37_io_dataRead)
  );
  Memory_108 spriteMemories_38 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_38_clock),
    .io_address(spriteMemories_38_io_address),
    .io_dataRead(spriteMemories_38_io_dataRead)
  );
  Memory_109 spriteMemories_39 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_39_clock),
    .io_address(spriteMemories_39_io_address),
    .io_dataRead(spriteMemories_39_io_dataRead)
  );
  Memory_110 spriteMemories_40 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_40_clock),
    .io_address(spriteMemories_40_io_address),
    .io_dataRead(spriteMemories_40_io_dataRead)
  );
  Memory_111 spriteMemories_41 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_41_clock),
    .io_address(spriteMemories_41_io_address),
    .io_dataRead(spriteMemories_41_io_dataRead)
  );
  Memory_112 spriteMemories_42 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_42_clock),
    .io_address(spriteMemories_42_io_address),
    .io_dataRead(spriteMemories_42_io_dataRead)
  );
  Memory_113 spriteMemories_43 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_43_clock),
    .io_address(spriteMemories_43_io_address),
    .io_dataRead(spriteMemories_43_io_dataRead)
  );
  Memory_114 spriteMemories_44 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_44_clock),
    .io_address(spriteMemories_44_io_address),
    .io_dataRead(spriteMemories_44_io_dataRead)
  );
  Memory_115 spriteMemories_45 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_45_clock),
    .io_address(spriteMemories_45_io_address),
    .io_dataRead(spriteMemories_45_io_dataRead)
  );
  Memory_116 spriteMemories_46 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_46_clock),
    .io_address(spriteMemories_46_io_address),
    .io_dataRead(spriteMemories_46_io_dataRead)
  );
  Memory_117 spriteMemories_47 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_47_clock),
    .io_address(spriteMemories_47_io_address),
    .io_dataRead(spriteMemories_47_io_dataRead)
  );
  Memory_118 spriteMemories_48 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_48_clock),
    .io_address(spriteMemories_48_io_address),
    .io_dataRead(spriteMemories_48_io_dataRead)
  );
  Memory_119 spriteMemories_49 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_49_clock),
    .io_address(spriteMemories_49_io_address),
    .io_dataRead(spriteMemories_49_io_dataRead)
  );
  Memory_120 spriteMemories_50 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_50_clock),
    .io_address(spriteMemories_50_io_address),
    .io_dataRead(spriteMemories_50_io_dataRead)
  );
  Memory_121 spriteMemories_51 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_51_clock),
    .io_address(spriteMemories_51_io_address),
    .io_dataRead(spriteMemories_51_io_dataRead)
  );
  Memory_122 spriteMemories_52 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_52_clock),
    .io_address(spriteMemories_52_io_address),
    .io_dataRead(spriteMemories_52_io_dataRead)
  );
  Memory_123 spriteMemories_53 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_53_clock),
    .io_address(spriteMemories_53_io_address),
    .io_dataRead(spriteMemories_53_io_dataRead)
  );
  Memory_124 spriteMemories_54 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_54_clock),
    .io_address(spriteMemories_54_io_address),
    .io_dataRead(spriteMemories_54_io_dataRead)
  );
  Memory_125 spriteMemories_55 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_55_clock),
    .io_address(spriteMemories_55_io_address),
    .io_dataRead(spriteMemories_55_io_dataRead)
  );
  Memory_126 spriteMemories_56 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_56_clock),
    .io_address(spriteMemories_56_io_address),
    .io_dataRead(spriteMemories_56_io_dataRead)
  );
  Memory_127 spriteMemories_57 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_57_clock),
    .io_address(spriteMemories_57_io_address),
    .io_dataRead(spriteMemories_57_io_dataRead)
  );
  Memory_128 spriteMemories_58 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_58_clock),
    .io_address(spriteMemories_58_io_address),
    .io_dataRead(spriteMemories_58_io_dataRead)
  );
  Memory_129 spriteMemories_59 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_59_clock),
    .io_address(spriteMemories_59_io_address),
    .io_dataRead(spriteMemories_59_io_dataRead)
  );
  Memory_130 spriteMemories_60 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_60_clock),
    .io_address(spriteMemories_60_io_address),
    .io_dataRead(spriteMemories_60_io_dataRead)
  );
  Memory_131 spriteMemories_61 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_61_clock),
    .io_address(spriteMemories_61_io_address),
    .io_dataRead(spriteMemories_61_io_dataRead)
  );
  Memory_132 spriteMemories_62 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_62_clock),
    .io_address(spriteMemories_62_io_address),
    .io_dataRead(spriteMemories_62_io_dataRead)
  );
  Memory_133 spriteMemories_63 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_63_clock),
    .io_address(spriteMemories_63_io_address),
    .io_dataRead(spriteMemories_63_io_dataRead)
  );
  Memory_134 spriteMemories_64 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_64_clock),
    .io_address(spriteMemories_64_io_address),
    .io_dataRead(spriteMemories_64_io_dataRead)
  );
  Memory_135 spriteMemories_65 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_65_clock),
    .io_address(spriteMemories_65_io_address),
    .io_dataRead(spriteMemories_65_io_dataRead)
  );
  Memory_136 spriteMemories_66 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_66_clock),
    .io_address(spriteMemories_66_io_address),
    .io_dataRead(spriteMemories_66_io_dataRead)
  );
  Memory_137 spriteMemories_67 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_67_clock),
    .io_address(spriteMemories_67_io_address),
    .io_dataRead(spriteMemories_67_io_dataRead)
  );
  Memory_138 spriteMemories_68 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_68_clock),
    .io_address(spriteMemories_68_io_address),
    .io_dataRead(spriteMemories_68_io_dataRead)
  );
  Memory_139 spriteMemories_69 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_69_clock),
    .io_address(spriteMemories_69_io_address),
    .io_dataRead(spriteMemories_69_io_dataRead)
  );
  Memory_140 spriteMemories_70 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_70_clock),
    .io_address(spriteMemories_70_io_address),
    .io_dataRead(spriteMemories_70_io_dataRead)
  );
  Memory_141 spriteMemories_71 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_71_clock),
    .io_address(spriteMemories_71_io_address),
    .io_dataRead(spriteMemories_71_io_dataRead)
  );
  Memory_142 spriteMemories_72 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_72_clock),
    .io_address(spriteMemories_72_io_address),
    .io_dataRead(spriteMemories_72_io_dataRead)
  );
  Memory_143 spriteMemories_73 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_73_clock),
    .io_address(spriteMemories_73_io_address),
    .io_dataRead(spriteMemories_73_io_dataRead)
  );
  Memory_144 spriteMemories_74 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_74_clock),
    .io_address(spriteMemories_74_io_address),
    .io_dataRead(spriteMemories_74_io_dataRead)
  );
  Memory_145 spriteMemories_75 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_75_clock),
    .io_address(spriteMemories_75_io_address),
    .io_dataRead(spriteMemories_75_io_dataRead)
  );
  Memory_146 spriteMemories_76 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_76_clock),
    .io_address(spriteMemories_76_io_address),
    .io_dataRead(spriteMemories_76_io_dataRead)
  );
  Memory_147 spriteMemories_77 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_77_clock),
    .io_address(spriteMemories_77_io_address),
    .io_dataRead(spriteMemories_77_io_dataRead)
  );
  Memory_148 spriteMemories_78 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_78_clock),
    .io_address(spriteMemories_78_io_address),
    .io_dataRead(spriteMemories_78_io_dataRead)
  );
  Memory_149 spriteMemories_79 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_79_clock),
    .io_address(spriteMemories_79_io_address),
    .io_dataRead(spriteMemories_79_io_dataRead)
  );
  Memory_150 spriteMemories_80 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_80_clock),
    .io_address(spriteMemories_80_io_address),
    .io_dataRead(spriteMemories_80_io_dataRead)
  );
  Memory_151 spriteMemories_81 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_81_clock),
    .io_address(spriteMemories_81_io_address),
    .io_dataRead(spriteMemories_81_io_dataRead)
  );
  Memory_152 spriteMemories_82 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_82_clock),
    .io_address(spriteMemories_82_io_address),
    .io_dataRead(spriteMemories_82_io_dataRead)
  );
  Memory_153 spriteMemories_83 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_83_clock),
    .io_address(spriteMemories_83_io_address),
    .io_dataRead(spriteMemories_83_io_dataRead)
  );
  Memory_154 spriteMemories_84 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_84_clock),
    .io_address(spriteMemories_84_io_address),
    .io_dataRead(spriteMemories_84_io_dataRead)
  );
  Memory_155 spriteMemories_85 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_85_clock),
    .io_address(spriteMemories_85_io_address),
    .io_dataRead(spriteMemories_85_io_dataRead)
  );
  Memory_156 spriteMemories_86 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_86_clock),
    .io_address(spriteMemories_86_io_address),
    .io_dataRead(spriteMemories_86_io_dataRead)
  );
  Memory_157 spriteMemories_87 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_87_clock),
    .io_address(spriteMemories_87_io_address),
    .io_dataRead(spriteMemories_87_io_dataRead)
  );
  Memory_158 spriteMemories_88 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_88_clock),
    .io_address(spriteMemories_88_io_address),
    .io_dataRead(spriteMemories_88_io_dataRead)
  );
  Memory_159 spriteMemories_89 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_89_clock),
    .io_address(spriteMemories_89_io_address),
    .io_dataRead(spriteMemories_89_io_dataRead)
  );
  Memory_160 spriteMemories_90 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_90_clock),
    .io_address(spriteMemories_90_io_address),
    .io_dataRead(spriteMemories_90_io_dataRead)
  );
  Memory_161 spriteMemories_91 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_91_clock),
    .io_address(spriteMemories_91_io_address),
    .io_dataRead(spriteMemories_91_io_dataRead)
  );
  Memory_162 spriteMemories_92 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_92_clock),
    .io_address(spriteMemories_92_io_address),
    .io_dataRead(spriteMemories_92_io_dataRead)
  );
  Memory_163 spriteMemories_93 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_93_clock),
    .io_address(spriteMemories_93_io_address),
    .io_dataRead(spriteMemories_93_io_dataRead)
  );
  Memory_164 spriteMemories_94 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_94_clock),
    .io_address(spriteMemories_94_io_address),
    .io_dataRead(spriteMemories_94_io_dataRead)
  );
  Memory_165 spriteMemories_95 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_95_clock),
    .io_address(spriteMemories_95_io_address),
    .io_dataRead(spriteMemories_95_io_dataRead)
  );
  Memory_166 spriteMemories_96 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_96_clock),
    .io_address(spriteMemories_96_io_address),
    .io_dataRead(spriteMemories_96_io_dataRead)
  );
  Memory_167 spriteMemories_97 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_97_clock),
    .io_address(spriteMemories_97_io_address),
    .io_dataRead(spriteMemories_97_io_dataRead)
  );
  Memory_168 spriteMemories_98 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_98_clock),
    .io_address(spriteMemories_98_io_address),
    .io_dataRead(spriteMemories_98_io_dataRead)
  );
  Memory_169 spriteMemories_99 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_99_clock),
    .io_address(spriteMemories_99_io_address),
    .io_dataRead(spriteMemories_99_io_dataRead)
  );
  Memory_170 spriteMemories_100 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_100_clock),
    .io_address(spriteMemories_100_io_address),
    .io_dataRead(spriteMemories_100_io_dataRead)
  );
  Memory_171 spriteMemories_101 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_101_clock),
    .io_address(spriteMemories_101_io_address),
    .io_dataRead(spriteMemories_101_io_dataRead)
  );
  Memory_172 spriteMemories_102 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_102_clock),
    .io_address(spriteMemories_102_io_address),
    .io_dataRead(spriteMemories_102_io_dataRead)
  );
  Memory_173 spriteMemories_103 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_103_clock),
    .io_address(spriteMemories_103_io_address),
    .io_dataRead(spriteMemories_103_io_dataRead)
  );
  Memory_174 spriteMemories_104 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_104_clock),
    .io_address(spriteMemories_104_io_address),
    .io_dataRead(spriteMemories_104_io_dataRead)
  );
  Memory_175 spriteMemories_105 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_105_clock),
    .io_address(spriteMemories_105_io_address),
    .io_dataRead(spriteMemories_105_io_dataRead)
  );
  Memory_176 spriteMemories_106 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_106_clock),
    .io_address(spriteMemories_106_io_address),
    .io_dataRead(spriteMemories_106_io_dataRead)
  );
  Memory_177 spriteMemories_107 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_107_clock),
    .io_address(spriteMemories_107_io_address),
    .io_dataRead(spriteMemories_107_io_dataRead)
  );
  Memory_178 spriteMemories_108 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_108_clock),
    .io_address(spriteMemories_108_io_address),
    .io_dataRead(spriteMemories_108_io_dataRead)
  );
  Memory_179 spriteMemories_109 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_109_clock),
    .io_address(spriteMemories_109_io_address),
    .io_dataRead(spriteMemories_109_io_dataRead)
  );
  Memory_180 spriteMemories_110 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_110_clock),
    .io_address(spriteMemories_110_io_address),
    .io_dataRead(spriteMemories_110_io_dataRead)
  );
  Memory_181 spriteMemories_111 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_111_clock),
    .io_address(spriteMemories_111_io_address),
    .io_dataRead(spriteMemories_111_io_dataRead)
  );
  Memory_182 spriteMemories_112 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_112_clock),
    .io_address(spriteMemories_112_io_address),
    .io_dataRead(spriteMemories_112_io_dataRead)
  );
  Memory_183 spriteMemories_113 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_113_clock),
    .io_address(spriteMemories_113_io_address),
    .io_dataRead(spriteMemories_113_io_dataRead)
  );
  Memory_184 spriteMemories_114 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_114_clock),
    .io_address(spriteMemories_114_io_address),
    .io_dataRead(spriteMemories_114_io_dataRead)
  );
  Memory_185 spriteMemories_115 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_115_clock),
    .io_address(spriteMemories_115_io_address),
    .io_dataRead(spriteMemories_115_io_dataRead)
  );
  Memory_186 spriteMemories_116 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_116_clock),
    .io_address(spriteMemories_116_io_address),
    .io_dataRead(spriteMemories_116_io_dataRead)
  );
  Memory_187 spriteMemories_117 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_117_clock),
    .io_address(spriteMemories_117_io_address),
    .io_dataRead(spriteMemories_117_io_dataRead)
  );
  Memory_188 spriteMemories_118 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_118_clock),
    .io_address(spriteMemories_118_io_address),
    .io_dataRead(spriteMemories_118_io_dataRead)
  );
  Memory_189 spriteMemories_119 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_119_clock),
    .io_address(spriteMemories_119_io_address),
    .io_dataRead(spriteMemories_119_io_dataRead)
  );
  Memory_190 spriteMemories_120 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_120_clock),
    .io_address(spriteMemories_120_io_address),
    .io_dataRead(spriteMemories_120_io_dataRead)
  );
  Memory_191 spriteMemories_121 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_121_clock),
    .io_address(spriteMemories_121_io_address),
    .io_dataRead(spriteMemories_121_io_dataRead)
  );
  Memory_192 spriteMemories_122 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_122_clock),
    .io_address(spriteMemories_122_io_address),
    .io_dataRead(spriteMemories_122_io_dataRead)
  );
  Memory_193 spriteMemories_123 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_123_clock),
    .io_address(spriteMemories_123_io_address),
    .io_dataRead(spriteMemories_123_io_dataRead)
  );
  Memory_194 spriteMemories_124 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_124_clock),
    .io_address(spriteMemories_124_io_address),
    .io_dataRead(spriteMemories_124_io_dataRead)
  );
  Memory_195 spriteMemories_125 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_125_clock),
    .io_address(spriteMemories_125_io_address),
    .io_dataRead(spriteMemories_125_io_dataRead)
  );
  Memory_196 spriteMemories_126 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_126_clock),
    .io_address(spriteMemories_126_io_address),
    .io_dataRead(spriteMemories_126_io_dataRead)
  );
  Memory_197 spriteMemories_127 ( // @[GraphicEngineVGA.scala 273:30]
    .clock(spriteMemories_127_clock),
    .io_address(spriteMemories_127_io_address),
    .io_dataRead(spriteMemories_127_io_dataRead)
  );
  MultiHotPriortyReductionTree multiHotPriortyReductionTree ( // @[GraphicEngineVGA.scala 306:44]
    .io_dataInput_0(multiHotPriortyReductionTree_io_dataInput_0),
    .io_dataInput_1(multiHotPriortyReductionTree_io_dataInput_1),
    .io_dataInput_2(multiHotPriortyReductionTree_io_dataInput_2),
    .io_dataInput_3(multiHotPriortyReductionTree_io_dataInput_3),
    .io_dataInput_4(multiHotPriortyReductionTree_io_dataInput_4),
    .io_dataInput_5(multiHotPriortyReductionTree_io_dataInput_5),
    .io_dataInput_6(multiHotPriortyReductionTree_io_dataInput_6),
    .io_dataInput_7(multiHotPriortyReductionTree_io_dataInput_7),
    .io_dataInput_8(multiHotPriortyReductionTree_io_dataInput_8),
    .io_dataInput_9(multiHotPriortyReductionTree_io_dataInput_9),
    .io_dataInput_10(multiHotPriortyReductionTree_io_dataInput_10),
    .io_dataInput_11(multiHotPriortyReductionTree_io_dataInput_11),
    .io_dataInput_12(multiHotPriortyReductionTree_io_dataInput_12),
    .io_dataInput_13(multiHotPriortyReductionTree_io_dataInput_13),
    .io_dataInput_14(multiHotPriortyReductionTree_io_dataInput_14),
    .io_dataInput_15(multiHotPriortyReductionTree_io_dataInput_15),
    .io_dataInput_16(multiHotPriortyReductionTree_io_dataInput_16),
    .io_dataInput_17(multiHotPriortyReductionTree_io_dataInput_17),
    .io_dataInput_18(multiHotPriortyReductionTree_io_dataInput_18),
    .io_dataInput_19(multiHotPriortyReductionTree_io_dataInput_19),
    .io_dataInput_20(multiHotPriortyReductionTree_io_dataInput_20),
    .io_dataInput_21(multiHotPriortyReductionTree_io_dataInput_21),
    .io_dataInput_22(multiHotPriortyReductionTree_io_dataInput_22),
    .io_dataInput_23(multiHotPriortyReductionTree_io_dataInput_23),
    .io_dataInput_24(multiHotPriortyReductionTree_io_dataInput_24),
    .io_dataInput_25(multiHotPriortyReductionTree_io_dataInput_25),
    .io_dataInput_26(multiHotPriortyReductionTree_io_dataInput_26),
    .io_dataInput_27(multiHotPriortyReductionTree_io_dataInput_27),
    .io_dataInput_28(multiHotPriortyReductionTree_io_dataInput_28),
    .io_dataInput_29(multiHotPriortyReductionTree_io_dataInput_29),
    .io_dataInput_30(multiHotPriortyReductionTree_io_dataInput_30),
    .io_dataInput_31(multiHotPriortyReductionTree_io_dataInput_31),
    .io_dataInput_32(multiHotPriortyReductionTree_io_dataInput_32),
    .io_dataInput_33(multiHotPriortyReductionTree_io_dataInput_33),
    .io_dataInput_34(multiHotPriortyReductionTree_io_dataInput_34),
    .io_dataInput_35(multiHotPriortyReductionTree_io_dataInput_35),
    .io_dataInput_36(multiHotPriortyReductionTree_io_dataInput_36),
    .io_dataInput_37(multiHotPriortyReductionTree_io_dataInput_37),
    .io_dataInput_38(multiHotPriortyReductionTree_io_dataInput_38),
    .io_dataInput_39(multiHotPriortyReductionTree_io_dataInput_39),
    .io_dataInput_40(multiHotPriortyReductionTree_io_dataInput_40),
    .io_dataInput_41(multiHotPriortyReductionTree_io_dataInput_41),
    .io_dataInput_42(multiHotPriortyReductionTree_io_dataInput_42),
    .io_dataInput_43(multiHotPriortyReductionTree_io_dataInput_43),
    .io_dataInput_44(multiHotPriortyReductionTree_io_dataInput_44),
    .io_dataInput_45(multiHotPriortyReductionTree_io_dataInput_45),
    .io_dataInput_46(multiHotPriortyReductionTree_io_dataInput_46),
    .io_dataInput_47(multiHotPriortyReductionTree_io_dataInput_47),
    .io_dataInput_48(multiHotPriortyReductionTree_io_dataInput_48),
    .io_dataInput_49(multiHotPriortyReductionTree_io_dataInput_49),
    .io_dataInput_50(multiHotPriortyReductionTree_io_dataInput_50),
    .io_dataInput_51(multiHotPriortyReductionTree_io_dataInput_51),
    .io_dataInput_52(multiHotPriortyReductionTree_io_dataInput_52),
    .io_dataInput_53(multiHotPriortyReductionTree_io_dataInput_53),
    .io_dataInput_54(multiHotPriortyReductionTree_io_dataInput_54),
    .io_dataInput_55(multiHotPriortyReductionTree_io_dataInput_55),
    .io_dataInput_56(multiHotPriortyReductionTree_io_dataInput_56),
    .io_dataInput_57(multiHotPriortyReductionTree_io_dataInput_57),
    .io_dataInput_58(multiHotPriortyReductionTree_io_dataInput_58),
    .io_dataInput_59(multiHotPriortyReductionTree_io_dataInput_59),
    .io_dataInput_60(multiHotPriortyReductionTree_io_dataInput_60),
    .io_dataInput_61(multiHotPriortyReductionTree_io_dataInput_61),
    .io_dataInput_62(multiHotPriortyReductionTree_io_dataInput_62),
    .io_dataInput_63(multiHotPriortyReductionTree_io_dataInput_63),
    .io_dataInput_64(multiHotPriortyReductionTree_io_dataInput_64),
    .io_dataInput_65(multiHotPriortyReductionTree_io_dataInput_65),
    .io_dataInput_66(multiHotPriortyReductionTree_io_dataInput_66),
    .io_dataInput_67(multiHotPriortyReductionTree_io_dataInput_67),
    .io_dataInput_68(multiHotPriortyReductionTree_io_dataInput_68),
    .io_dataInput_69(multiHotPriortyReductionTree_io_dataInput_69),
    .io_dataInput_70(multiHotPriortyReductionTree_io_dataInput_70),
    .io_dataInput_71(multiHotPriortyReductionTree_io_dataInput_71),
    .io_dataInput_72(multiHotPriortyReductionTree_io_dataInput_72),
    .io_dataInput_73(multiHotPriortyReductionTree_io_dataInput_73),
    .io_dataInput_74(multiHotPriortyReductionTree_io_dataInput_74),
    .io_dataInput_75(multiHotPriortyReductionTree_io_dataInput_75),
    .io_dataInput_76(multiHotPriortyReductionTree_io_dataInput_76),
    .io_dataInput_77(multiHotPriortyReductionTree_io_dataInput_77),
    .io_dataInput_78(multiHotPriortyReductionTree_io_dataInput_78),
    .io_dataInput_79(multiHotPriortyReductionTree_io_dataInput_79),
    .io_dataInput_80(multiHotPriortyReductionTree_io_dataInput_80),
    .io_dataInput_81(multiHotPriortyReductionTree_io_dataInput_81),
    .io_dataInput_82(multiHotPriortyReductionTree_io_dataInput_82),
    .io_dataInput_83(multiHotPriortyReductionTree_io_dataInput_83),
    .io_dataInput_84(multiHotPriortyReductionTree_io_dataInput_84),
    .io_dataInput_85(multiHotPriortyReductionTree_io_dataInput_85),
    .io_dataInput_86(multiHotPriortyReductionTree_io_dataInput_86),
    .io_dataInput_87(multiHotPriortyReductionTree_io_dataInput_87),
    .io_dataInput_88(multiHotPriortyReductionTree_io_dataInput_88),
    .io_dataInput_89(multiHotPriortyReductionTree_io_dataInput_89),
    .io_dataInput_90(multiHotPriortyReductionTree_io_dataInput_90),
    .io_dataInput_91(multiHotPriortyReductionTree_io_dataInput_91),
    .io_dataInput_92(multiHotPriortyReductionTree_io_dataInput_92),
    .io_dataInput_93(multiHotPriortyReductionTree_io_dataInput_93),
    .io_dataInput_94(multiHotPriortyReductionTree_io_dataInput_94),
    .io_dataInput_95(multiHotPriortyReductionTree_io_dataInput_95),
    .io_dataInput_96(multiHotPriortyReductionTree_io_dataInput_96),
    .io_dataInput_97(multiHotPriortyReductionTree_io_dataInput_97),
    .io_dataInput_98(multiHotPriortyReductionTree_io_dataInput_98),
    .io_dataInput_99(multiHotPriortyReductionTree_io_dataInput_99),
    .io_dataInput_100(multiHotPriortyReductionTree_io_dataInput_100),
    .io_dataInput_101(multiHotPriortyReductionTree_io_dataInput_101),
    .io_dataInput_102(multiHotPriortyReductionTree_io_dataInput_102),
    .io_dataInput_103(multiHotPriortyReductionTree_io_dataInput_103),
    .io_dataInput_104(multiHotPriortyReductionTree_io_dataInput_104),
    .io_dataInput_105(multiHotPriortyReductionTree_io_dataInput_105),
    .io_dataInput_106(multiHotPriortyReductionTree_io_dataInput_106),
    .io_dataInput_107(multiHotPriortyReductionTree_io_dataInput_107),
    .io_dataInput_108(multiHotPriortyReductionTree_io_dataInput_108),
    .io_dataInput_109(multiHotPriortyReductionTree_io_dataInput_109),
    .io_dataInput_110(multiHotPriortyReductionTree_io_dataInput_110),
    .io_dataInput_111(multiHotPriortyReductionTree_io_dataInput_111),
    .io_dataInput_112(multiHotPriortyReductionTree_io_dataInput_112),
    .io_dataInput_113(multiHotPriortyReductionTree_io_dataInput_113),
    .io_dataInput_114(multiHotPriortyReductionTree_io_dataInput_114),
    .io_dataInput_115(multiHotPriortyReductionTree_io_dataInput_115),
    .io_dataInput_116(multiHotPriortyReductionTree_io_dataInput_116),
    .io_dataInput_117(multiHotPriortyReductionTree_io_dataInput_117),
    .io_dataInput_118(multiHotPriortyReductionTree_io_dataInput_118),
    .io_dataInput_119(multiHotPriortyReductionTree_io_dataInput_119),
    .io_dataInput_120(multiHotPriortyReductionTree_io_dataInput_120),
    .io_dataInput_121(multiHotPriortyReductionTree_io_dataInput_121),
    .io_dataInput_122(multiHotPriortyReductionTree_io_dataInput_122),
    .io_dataInput_123(multiHotPriortyReductionTree_io_dataInput_123),
    .io_dataInput_124(multiHotPriortyReductionTree_io_dataInput_124),
    .io_dataInput_125(multiHotPriortyReductionTree_io_dataInput_125),
    .io_dataInput_126(multiHotPriortyReductionTree_io_dataInput_126),
    .io_dataInput_127(multiHotPriortyReductionTree_io_dataInput_127),
    .io_selectInput_0(multiHotPriortyReductionTree_io_selectInput_0),
    .io_selectInput_1(multiHotPriortyReductionTree_io_selectInput_1),
    .io_selectInput_2(multiHotPriortyReductionTree_io_selectInput_2),
    .io_selectInput_3(multiHotPriortyReductionTree_io_selectInput_3),
    .io_selectInput_4(multiHotPriortyReductionTree_io_selectInput_4),
    .io_selectInput_5(multiHotPriortyReductionTree_io_selectInput_5),
    .io_selectInput_6(multiHotPriortyReductionTree_io_selectInput_6),
    .io_selectInput_7(multiHotPriortyReductionTree_io_selectInput_7),
    .io_selectInput_8(multiHotPriortyReductionTree_io_selectInput_8),
    .io_selectInput_9(multiHotPriortyReductionTree_io_selectInput_9),
    .io_selectInput_10(multiHotPriortyReductionTree_io_selectInput_10),
    .io_selectInput_11(multiHotPriortyReductionTree_io_selectInput_11),
    .io_selectInput_12(multiHotPriortyReductionTree_io_selectInput_12),
    .io_selectInput_13(multiHotPriortyReductionTree_io_selectInput_13),
    .io_selectInput_14(multiHotPriortyReductionTree_io_selectInput_14),
    .io_selectInput_15(multiHotPriortyReductionTree_io_selectInput_15),
    .io_selectInput_16(multiHotPriortyReductionTree_io_selectInput_16),
    .io_selectInput_17(multiHotPriortyReductionTree_io_selectInput_17),
    .io_selectInput_18(multiHotPriortyReductionTree_io_selectInput_18),
    .io_selectInput_19(multiHotPriortyReductionTree_io_selectInput_19),
    .io_selectInput_20(multiHotPriortyReductionTree_io_selectInput_20),
    .io_selectInput_21(multiHotPriortyReductionTree_io_selectInput_21),
    .io_selectInput_22(multiHotPriortyReductionTree_io_selectInput_22),
    .io_selectInput_23(multiHotPriortyReductionTree_io_selectInput_23),
    .io_selectInput_24(multiHotPriortyReductionTree_io_selectInput_24),
    .io_selectInput_25(multiHotPriortyReductionTree_io_selectInput_25),
    .io_selectInput_26(multiHotPriortyReductionTree_io_selectInput_26),
    .io_selectInput_27(multiHotPriortyReductionTree_io_selectInput_27),
    .io_selectInput_28(multiHotPriortyReductionTree_io_selectInput_28),
    .io_selectInput_29(multiHotPriortyReductionTree_io_selectInput_29),
    .io_selectInput_30(multiHotPriortyReductionTree_io_selectInput_30),
    .io_selectInput_31(multiHotPriortyReductionTree_io_selectInput_31),
    .io_selectInput_32(multiHotPriortyReductionTree_io_selectInput_32),
    .io_selectInput_33(multiHotPriortyReductionTree_io_selectInput_33),
    .io_selectInput_34(multiHotPriortyReductionTree_io_selectInput_34),
    .io_selectInput_35(multiHotPriortyReductionTree_io_selectInput_35),
    .io_selectInput_36(multiHotPriortyReductionTree_io_selectInput_36),
    .io_selectInput_37(multiHotPriortyReductionTree_io_selectInput_37),
    .io_selectInput_38(multiHotPriortyReductionTree_io_selectInput_38),
    .io_selectInput_39(multiHotPriortyReductionTree_io_selectInput_39),
    .io_selectInput_40(multiHotPriortyReductionTree_io_selectInput_40),
    .io_selectInput_41(multiHotPriortyReductionTree_io_selectInput_41),
    .io_selectInput_42(multiHotPriortyReductionTree_io_selectInput_42),
    .io_selectInput_43(multiHotPriortyReductionTree_io_selectInput_43),
    .io_selectInput_44(multiHotPriortyReductionTree_io_selectInput_44),
    .io_selectInput_45(multiHotPriortyReductionTree_io_selectInput_45),
    .io_selectInput_46(multiHotPriortyReductionTree_io_selectInput_46),
    .io_selectInput_47(multiHotPriortyReductionTree_io_selectInput_47),
    .io_selectInput_48(multiHotPriortyReductionTree_io_selectInput_48),
    .io_selectInput_49(multiHotPriortyReductionTree_io_selectInput_49),
    .io_selectInput_50(multiHotPriortyReductionTree_io_selectInput_50),
    .io_selectInput_51(multiHotPriortyReductionTree_io_selectInput_51),
    .io_selectInput_52(multiHotPriortyReductionTree_io_selectInput_52),
    .io_selectInput_53(multiHotPriortyReductionTree_io_selectInput_53),
    .io_selectInput_54(multiHotPriortyReductionTree_io_selectInput_54),
    .io_selectInput_55(multiHotPriortyReductionTree_io_selectInput_55),
    .io_selectInput_56(multiHotPriortyReductionTree_io_selectInput_56),
    .io_selectInput_57(multiHotPriortyReductionTree_io_selectInput_57),
    .io_selectInput_58(multiHotPriortyReductionTree_io_selectInput_58),
    .io_selectInput_59(multiHotPriortyReductionTree_io_selectInput_59),
    .io_selectInput_60(multiHotPriortyReductionTree_io_selectInput_60),
    .io_selectInput_61(multiHotPriortyReductionTree_io_selectInput_61),
    .io_selectInput_62(multiHotPriortyReductionTree_io_selectInput_62),
    .io_selectInput_63(multiHotPriortyReductionTree_io_selectInput_63),
    .io_selectInput_64(multiHotPriortyReductionTree_io_selectInput_64),
    .io_selectInput_65(multiHotPriortyReductionTree_io_selectInput_65),
    .io_selectInput_66(multiHotPriortyReductionTree_io_selectInput_66),
    .io_selectInput_67(multiHotPriortyReductionTree_io_selectInput_67),
    .io_selectInput_68(multiHotPriortyReductionTree_io_selectInput_68),
    .io_selectInput_69(multiHotPriortyReductionTree_io_selectInput_69),
    .io_selectInput_70(multiHotPriortyReductionTree_io_selectInput_70),
    .io_selectInput_71(multiHotPriortyReductionTree_io_selectInput_71),
    .io_selectInput_72(multiHotPriortyReductionTree_io_selectInput_72),
    .io_selectInput_73(multiHotPriortyReductionTree_io_selectInput_73),
    .io_selectInput_74(multiHotPriortyReductionTree_io_selectInput_74),
    .io_selectInput_75(multiHotPriortyReductionTree_io_selectInput_75),
    .io_selectInput_76(multiHotPriortyReductionTree_io_selectInput_76),
    .io_selectInput_77(multiHotPriortyReductionTree_io_selectInput_77),
    .io_selectInput_78(multiHotPriortyReductionTree_io_selectInput_78),
    .io_selectInput_79(multiHotPriortyReductionTree_io_selectInput_79),
    .io_selectInput_80(multiHotPriortyReductionTree_io_selectInput_80),
    .io_selectInput_81(multiHotPriortyReductionTree_io_selectInput_81),
    .io_selectInput_82(multiHotPriortyReductionTree_io_selectInput_82),
    .io_selectInput_83(multiHotPriortyReductionTree_io_selectInput_83),
    .io_selectInput_84(multiHotPriortyReductionTree_io_selectInput_84),
    .io_selectInput_85(multiHotPriortyReductionTree_io_selectInput_85),
    .io_selectInput_86(multiHotPriortyReductionTree_io_selectInput_86),
    .io_selectInput_87(multiHotPriortyReductionTree_io_selectInput_87),
    .io_selectInput_88(multiHotPriortyReductionTree_io_selectInput_88),
    .io_selectInput_89(multiHotPriortyReductionTree_io_selectInput_89),
    .io_selectInput_90(multiHotPriortyReductionTree_io_selectInput_90),
    .io_selectInput_91(multiHotPriortyReductionTree_io_selectInput_91),
    .io_selectInput_92(multiHotPriortyReductionTree_io_selectInput_92),
    .io_selectInput_93(multiHotPriortyReductionTree_io_selectInput_93),
    .io_selectInput_94(multiHotPriortyReductionTree_io_selectInput_94),
    .io_selectInput_95(multiHotPriortyReductionTree_io_selectInput_95),
    .io_selectInput_96(multiHotPriortyReductionTree_io_selectInput_96),
    .io_selectInput_97(multiHotPriortyReductionTree_io_selectInput_97),
    .io_selectInput_98(multiHotPriortyReductionTree_io_selectInput_98),
    .io_selectInput_99(multiHotPriortyReductionTree_io_selectInput_99),
    .io_selectInput_100(multiHotPriortyReductionTree_io_selectInput_100),
    .io_selectInput_101(multiHotPriortyReductionTree_io_selectInput_101),
    .io_selectInput_102(multiHotPriortyReductionTree_io_selectInput_102),
    .io_selectInput_103(multiHotPriortyReductionTree_io_selectInput_103),
    .io_selectInput_104(multiHotPriortyReductionTree_io_selectInput_104),
    .io_selectInput_105(multiHotPriortyReductionTree_io_selectInput_105),
    .io_selectInput_106(multiHotPriortyReductionTree_io_selectInput_106),
    .io_selectInput_107(multiHotPriortyReductionTree_io_selectInput_107),
    .io_selectInput_108(multiHotPriortyReductionTree_io_selectInput_108),
    .io_selectInput_109(multiHotPriortyReductionTree_io_selectInput_109),
    .io_selectInput_110(multiHotPriortyReductionTree_io_selectInput_110),
    .io_selectInput_111(multiHotPriortyReductionTree_io_selectInput_111),
    .io_selectInput_112(multiHotPriortyReductionTree_io_selectInput_112),
    .io_selectInput_113(multiHotPriortyReductionTree_io_selectInput_113),
    .io_selectInput_114(multiHotPriortyReductionTree_io_selectInput_114),
    .io_selectInput_115(multiHotPriortyReductionTree_io_selectInput_115),
    .io_selectInput_116(multiHotPriortyReductionTree_io_selectInput_116),
    .io_selectInput_117(multiHotPriortyReductionTree_io_selectInput_117),
    .io_selectInput_118(multiHotPriortyReductionTree_io_selectInput_118),
    .io_selectInput_119(multiHotPriortyReductionTree_io_selectInput_119),
    .io_selectInput_120(multiHotPriortyReductionTree_io_selectInput_120),
    .io_selectInput_121(multiHotPriortyReductionTree_io_selectInput_121),
    .io_selectInput_122(multiHotPriortyReductionTree_io_selectInput_122),
    .io_selectInput_123(multiHotPriortyReductionTree_io_selectInput_123),
    .io_selectInput_124(multiHotPriortyReductionTree_io_selectInput_124),
    .io_selectInput_125(multiHotPriortyReductionTree_io_selectInput_125),
    .io_selectInput_126(multiHotPriortyReductionTree_io_selectInput_126),
    .io_selectInput_127(multiHotPriortyReductionTree_io_selectInput_127),
    .io_dataOutput(multiHotPriortyReductionTree_io_dataOutput),
    .io_selectOutput(multiHotPriortyReductionTree_io_selectOutput)
  );
  assign io_newFrame = run & _GEN_8; // @[GraphicEngineVGA.scala 67:15 GraphicEngineVGA.scala 76:23]
  assign io_missingFrameError = missingFrameErrorReg; // @[GraphicEngineVGA.scala 125:24]
  assign io_backBufferWriteError = backBufferWriteErrorReg; // @[GraphicEngineVGA.scala 126:27]
  assign io_viewBoxOutOfRangeError = viewBoxOutOfRangeErrorReg; // @[GraphicEngineVGA.scala 127:29]
  assign io_vgaRed = _T_4655; // @[GraphicEngineVGA.scala 321:13]
  assign io_vgaBlue = _T_4657; // @[GraphicEngineVGA.scala 323:14]
  assign io_vgaGreen = _T_4656; // @[GraphicEngineVGA.scala 322:15]
  assign io_Hsync = _T_14_0; // @[GraphicEngineVGA.scala 90:12]
  assign io_Vsync = _T_16_0; // @[GraphicEngineVGA.scala 91:12]
  assign backTileMemories_0_0_clock = clock;
  assign backTileMemories_0_0_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_1_clock = clock;
  assign backTileMemories_0_1_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_2_clock = clock;
  assign backTileMemories_0_2_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_3_clock = clock;
  assign backTileMemories_0_3_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_4_clock = clock;
  assign backTileMemories_0_4_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_5_clock = clock;
  assign backTileMemories_0_5_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_6_clock = clock;
  assign backTileMemories_0_6_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_7_clock = clock;
  assign backTileMemories_0_7_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_8_clock = clock;
  assign backTileMemories_0_8_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_9_clock = clock;
  assign backTileMemories_0_9_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_10_clock = clock;
  assign backTileMemories_0_10_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_11_clock = clock;
  assign backTileMemories_0_11_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_12_clock = clock;
  assign backTileMemories_0_12_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_13_clock = clock;
  assign backTileMemories_0_13_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_14_clock = clock;
  assign backTileMemories_0_14_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_15_clock = clock;
  assign backTileMemories_0_15_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_16_clock = clock;
  assign backTileMemories_0_16_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_17_clock = clock;
  assign backTileMemories_0_17_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_18_clock = clock;
  assign backTileMemories_0_18_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_19_clock = clock;
  assign backTileMemories_0_19_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_20_clock = clock;
  assign backTileMemories_0_20_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_21_clock = clock;
  assign backTileMemories_0_21_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_22_clock = clock;
  assign backTileMemories_0_22_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_23_clock = clock;
  assign backTileMemories_0_23_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_24_clock = clock;
  assign backTileMemories_0_24_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_25_clock = clock;
  assign backTileMemories_0_25_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_26_clock = clock;
  assign backTileMemories_0_26_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_27_clock = clock;
  assign backTileMemories_0_27_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_28_clock = clock;
  assign backTileMemories_0_28_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_29_clock = clock;
  assign backTileMemories_0_29_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_30_clock = clock;
  assign backTileMemories_0_30_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_0_31_clock = clock;
  assign backTileMemories_0_31_io_address = _T_48[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_0_clock = clock;
  assign backTileMemories_1_0_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_1_clock = clock;
  assign backTileMemories_1_1_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_2_clock = clock;
  assign backTileMemories_1_2_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_3_clock = clock;
  assign backTileMemories_1_3_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_4_clock = clock;
  assign backTileMemories_1_4_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_5_clock = clock;
  assign backTileMemories_1_5_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_6_clock = clock;
  assign backTileMemories_1_6_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_7_clock = clock;
  assign backTileMemories_1_7_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_8_clock = clock;
  assign backTileMemories_1_8_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_9_clock = clock;
  assign backTileMemories_1_9_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_10_clock = clock;
  assign backTileMemories_1_10_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_11_clock = clock;
  assign backTileMemories_1_11_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_12_clock = clock;
  assign backTileMemories_1_12_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_13_clock = clock;
  assign backTileMemories_1_13_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_14_clock = clock;
  assign backTileMemories_1_14_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_15_clock = clock;
  assign backTileMemories_1_15_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_16_clock = clock;
  assign backTileMemories_1_16_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_17_clock = clock;
  assign backTileMemories_1_17_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_18_clock = clock;
  assign backTileMemories_1_18_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_19_clock = clock;
  assign backTileMemories_1_19_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_20_clock = clock;
  assign backTileMemories_1_20_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_21_clock = clock;
  assign backTileMemories_1_21_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_22_clock = clock;
  assign backTileMemories_1_22_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_23_clock = clock;
  assign backTileMemories_1_23_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_24_clock = clock;
  assign backTileMemories_1_24_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_25_clock = clock;
  assign backTileMemories_1_25_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_26_clock = clock;
  assign backTileMemories_1_26_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_27_clock = clock;
  assign backTileMemories_1_27_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_28_clock = clock;
  assign backTileMemories_1_28_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_29_clock = clock;
  assign backTileMemories_1_29_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_30_clock = clock;
  assign backTileMemories_1_30_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backTileMemories_1_31_clock = clock;
  assign backTileMemories_1_31_io_address = _T_208[9:0]; // @[GraphicEngineVGA.scala 175:39]
  assign backBufferMemories_0_clock = clock;
  assign backBufferMemories_0_io_address = _T_390[10:0]; // @[GraphicEngineVGA.scala 245:36]
  assign backBufferMemories_0_io_writeEnable = copyEnabledReg; // @[GraphicEngineVGA.scala 247:40]
  assign backBufferMemories_0_io_dataWrite = backBufferShadowMemories_0_io_dataRead; // @[GraphicEngineVGA.scala 248:38]
  assign backBufferMemories_1_clock = clock;
  assign backBufferMemories_1_io_address = _T_410[10:0]; // @[GraphicEngineVGA.scala 245:36]
  assign backBufferMemories_1_io_writeEnable = copyEnabledReg; // @[GraphicEngineVGA.scala 247:40]
  assign backBufferMemories_1_io_dataWrite = backBufferShadowMemories_1_io_dataRead; // @[GraphicEngineVGA.scala 248:38]
  assign backBufferShadowMemories_0_clock = clock;
  assign backBufferShadowMemories_0_io_address = restoreEnabled ? _T_373 : _T_376; // @[GraphicEngineVGA.scala 240:42]
  assign backBufferShadowMemories_0_io_writeEnable = restoreEnabled ? _T_378 : _T_380; // @[GraphicEngineVGA.scala 242:46]
  assign backBufferShadowMemories_0_io_dataWrite = restoreEnabled ? backBufferRestoreMemories_0_io_dataRead : _T_382; // @[GraphicEngineVGA.scala 243:44]
  assign backBufferShadowMemories_1_clock = clock;
  assign backBufferShadowMemories_1_io_address = restoreEnabled ? _T_393 : _T_396; // @[GraphicEngineVGA.scala 240:42]
  assign backBufferShadowMemories_1_io_writeEnable = restoreEnabled ? _T_398 : _T_400; // @[GraphicEngineVGA.scala 242:46]
  assign backBufferShadowMemories_1_io_dataWrite = restoreEnabled ? backBufferRestoreMemories_1_io_dataRead : _T_402; // @[GraphicEngineVGA.scala 243:44]
  assign backBufferRestoreMemories_0_clock = clock;
  assign backBufferRestoreMemories_0_io_address = backMemoryRestoreCounter[10:0]; // @[GraphicEngineVGA.scala 235:43]
  assign backBufferRestoreMemories_1_clock = clock;
  assign backBufferRestoreMemories_1_io_address = backMemoryRestoreCounter[10:0]; // @[GraphicEngineVGA.scala 235:43]
  assign spriteMemories_0_clock = clock;
  assign spriteMemories_0_io_address = _T_2860[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_1_clock = clock;
  assign spriteMemories_1_io_address = _T_2865[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_2_clock = clock;
  assign spriteMemories_2_io_address = _T_2870[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_3_clock = clock;
  assign spriteMemories_3_io_address = _T_2875[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_4_clock = clock;
  assign spriteMemories_4_io_address = _T_2880[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_5_clock = clock;
  assign spriteMemories_5_io_address = _T_2885[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_6_clock = clock;
  assign spriteMemories_6_io_address = _T_2890[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_7_clock = clock;
  assign spriteMemories_7_io_address = _T_2895[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_8_clock = clock;
  assign spriteMemories_8_io_address = _T_2900[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_9_clock = clock;
  assign spriteMemories_9_io_address = _T_2905[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_10_clock = clock;
  assign spriteMemories_10_io_address = _T_2910[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_11_clock = clock;
  assign spriteMemories_11_io_address = _T_2915[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_12_clock = clock;
  assign spriteMemories_12_io_address = _T_2920[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_13_clock = clock;
  assign spriteMemories_13_io_address = _T_2925[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_14_clock = clock;
  assign spriteMemories_14_io_address = _T_2930[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_15_clock = clock;
  assign spriteMemories_15_io_address = _T_2935[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_16_clock = clock;
  assign spriteMemories_16_io_address = _T_2940[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_17_clock = clock;
  assign spriteMemories_17_io_address = _T_2945[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_18_clock = clock;
  assign spriteMemories_18_io_address = _T_2950[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_19_clock = clock;
  assign spriteMemories_19_io_address = _T_2955[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_20_clock = clock;
  assign spriteMemories_20_io_address = _T_2960[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_21_clock = clock;
  assign spriteMemories_21_io_address = _T_2965[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_22_clock = clock;
  assign spriteMemories_22_io_address = _T_2970[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_23_clock = clock;
  assign spriteMemories_23_io_address = _T_2975[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_24_clock = clock;
  assign spriteMemories_24_io_address = _T_2980[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_25_clock = clock;
  assign spriteMemories_25_io_address = _T_2985[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_26_clock = clock;
  assign spriteMemories_26_io_address = _T_2990[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_27_clock = clock;
  assign spriteMemories_27_io_address = _T_2995[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_28_clock = clock;
  assign spriteMemories_28_io_address = _T_3000[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_29_clock = clock;
  assign spriteMemories_29_io_address = _T_3005[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_30_clock = clock;
  assign spriteMemories_30_io_address = _T_3010[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_31_clock = clock;
  assign spriteMemories_31_io_address = _T_3015[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_32_clock = clock;
  assign spriteMemories_32_io_address = _T_3020[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_33_clock = clock;
  assign spriteMemories_33_io_address = _T_3025[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_34_clock = clock;
  assign spriteMemories_34_io_address = _T_3030[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_35_clock = clock;
  assign spriteMemories_35_io_address = _T_3035[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_36_clock = clock;
  assign spriteMemories_36_io_address = _T_3040[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_37_clock = clock;
  assign spriteMemories_37_io_address = _T_3045[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_38_clock = clock;
  assign spriteMemories_38_io_address = _T_3050[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_39_clock = clock;
  assign spriteMemories_39_io_address = _T_3055[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_40_clock = clock;
  assign spriteMemories_40_io_address = _T_3060[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_41_clock = clock;
  assign spriteMemories_41_io_address = _T_3065[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_42_clock = clock;
  assign spriteMemories_42_io_address = _T_3070[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_43_clock = clock;
  assign spriteMemories_43_io_address = _T_3075[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_44_clock = clock;
  assign spriteMemories_44_io_address = _T_3080[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_45_clock = clock;
  assign spriteMemories_45_io_address = _T_3085[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_46_clock = clock;
  assign spriteMemories_46_io_address = _T_3090[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_47_clock = clock;
  assign spriteMemories_47_io_address = _T_3095[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_48_clock = clock;
  assign spriteMemories_48_io_address = _T_3100[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_49_clock = clock;
  assign spriteMemories_49_io_address = _T_3105[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_50_clock = clock;
  assign spriteMemories_50_io_address = _T_3110[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_51_clock = clock;
  assign spriteMemories_51_io_address = _T_3115[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_52_clock = clock;
  assign spriteMemories_52_io_address = _T_3120[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_53_clock = clock;
  assign spriteMemories_53_io_address = _T_3125[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_54_clock = clock;
  assign spriteMemories_54_io_address = _T_3130[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_55_clock = clock;
  assign spriteMemories_55_io_address = _T_3135[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_56_clock = clock;
  assign spriteMemories_56_io_address = _T_3140[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_57_clock = clock;
  assign spriteMemories_57_io_address = _T_3145[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_58_clock = clock;
  assign spriteMemories_58_io_address = _T_3150[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_59_clock = clock;
  assign spriteMemories_59_io_address = _T_3155[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_60_clock = clock;
  assign spriteMemories_60_io_address = _T_3160[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_61_clock = clock;
  assign spriteMemories_61_io_address = _T_3165[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_62_clock = clock;
  assign spriteMemories_62_io_address = _T_3170[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_63_clock = clock;
  assign spriteMemories_63_io_address = _T_3175[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_64_clock = clock;
  assign spriteMemories_64_io_address = _T_3180[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_65_clock = clock;
  assign spriteMemories_65_io_address = _T_3185[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_66_clock = clock;
  assign spriteMemories_66_io_address = _T_3190[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_67_clock = clock;
  assign spriteMemories_67_io_address = _T_3195[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_68_clock = clock;
  assign spriteMemories_68_io_address = _T_3200[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_69_clock = clock;
  assign spriteMemories_69_io_address = _T_3205[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_70_clock = clock;
  assign spriteMemories_70_io_address = _T_3210[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_71_clock = clock;
  assign spriteMemories_71_io_address = _T_3215[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_72_clock = clock;
  assign spriteMemories_72_io_address = _T_3220[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_73_clock = clock;
  assign spriteMemories_73_io_address = _T_3225[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_74_clock = clock;
  assign spriteMemories_74_io_address = _T_3230[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_75_clock = clock;
  assign spriteMemories_75_io_address = _T_3235[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_76_clock = clock;
  assign spriteMemories_76_io_address = _T_3240[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_77_clock = clock;
  assign spriteMemories_77_io_address = _T_3245[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_78_clock = clock;
  assign spriteMemories_78_io_address = _T_3250[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_79_clock = clock;
  assign spriteMemories_79_io_address = _T_3255[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_80_clock = clock;
  assign spriteMemories_80_io_address = _T_3260[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_81_clock = clock;
  assign spriteMemories_81_io_address = _T_3265[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_82_clock = clock;
  assign spriteMemories_82_io_address = _T_3270[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_83_clock = clock;
  assign spriteMemories_83_io_address = _T_3275[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_84_clock = clock;
  assign spriteMemories_84_io_address = _T_3280[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_85_clock = clock;
  assign spriteMemories_85_io_address = _T_3285[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_86_clock = clock;
  assign spriteMemories_86_io_address = _T_3290[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_87_clock = clock;
  assign spriteMemories_87_io_address = _T_3295[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_88_clock = clock;
  assign spriteMemories_88_io_address = _T_3300[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_89_clock = clock;
  assign spriteMemories_89_io_address = _T_3305[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_90_clock = clock;
  assign spriteMemories_90_io_address = _T_3310[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_91_clock = clock;
  assign spriteMemories_91_io_address = _T_3315[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_92_clock = clock;
  assign spriteMemories_92_io_address = _T_3320[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_93_clock = clock;
  assign spriteMemories_93_io_address = _T_3325[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_94_clock = clock;
  assign spriteMemories_94_io_address = _T_3330[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_95_clock = clock;
  assign spriteMemories_95_io_address = _T_3335[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_96_clock = clock;
  assign spriteMemories_96_io_address = _T_3340[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_97_clock = clock;
  assign spriteMemories_97_io_address = _T_3345[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_98_clock = clock;
  assign spriteMemories_98_io_address = _T_3350[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_99_clock = clock;
  assign spriteMemories_99_io_address = _T_3355[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_100_clock = clock;
  assign spriteMemories_100_io_address = _T_3360[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_101_clock = clock;
  assign spriteMemories_101_io_address = _T_3365[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_102_clock = clock;
  assign spriteMemories_102_io_address = _T_3370[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_103_clock = clock;
  assign spriteMemories_103_io_address = _T_3375[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_104_clock = clock;
  assign spriteMemories_104_io_address = _T_3380[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_105_clock = clock;
  assign spriteMemories_105_io_address = _T_3385[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_106_clock = clock;
  assign spriteMemories_106_io_address = _T_3390[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_107_clock = clock;
  assign spriteMemories_107_io_address = _T_3395[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_108_clock = clock;
  assign spriteMemories_108_io_address = _T_3400[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_109_clock = clock;
  assign spriteMemories_109_io_address = _T_3405[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_110_clock = clock;
  assign spriteMemories_110_io_address = _T_3410[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_111_clock = clock;
  assign spriteMemories_111_io_address = _T_3415[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_112_clock = clock;
  assign spriteMemories_112_io_address = _T_3420[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_113_clock = clock;
  assign spriteMemories_113_io_address = _T_3425[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_114_clock = clock;
  assign spriteMemories_114_io_address = _T_3430[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_115_clock = clock;
  assign spriteMemories_115_io_address = _T_3435[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_116_clock = clock;
  assign spriteMemories_116_io_address = _T_3440[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_117_clock = clock;
  assign spriteMemories_117_io_address = _T_3445[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_118_clock = clock;
  assign spriteMemories_118_io_address = _T_3450[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_119_clock = clock;
  assign spriteMemories_119_io_address = _T_3455[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_120_clock = clock;
  assign spriteMemories_120_io_address = _T_3460[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_121_clock = clock;
  assign spriteMemories_121_io_address = _T_3465[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_122_clock = clock;
  assign spriteMemories_122_io_address = _T_3470[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_123_clock = clock;
  assign spriteMemories_123_io_address = _T_3475[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_124_clock = clock;
  assign spriteMemories_124_io_address = _T_3480[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_125_clock = clock;
  assign spriteMemories_125_io_address = _T_3485[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_126_clock = clock;
  assign spriteMemories_126_io_address = _T_3490[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign spriteMemories_127_clock = clock;
  assign spriteMemories_127_io_address = _T_3495[9:0]; // @[GraphicEngineVGA.scala 301:34]
  assign multiHotPriortyReductionTree_io_dataInput_0 = _T_3497; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_1 = _T_3506; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_2 = _T_3515; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_3 = _T_3524; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_4 = _T_3533; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_5 = _T_3542; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_6 = _T_3551; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_7 = _T_3560; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_8 = _T_3569; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_9 = _T_3578; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_10 = _T_3587; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_11 = _T_3596; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_12 = _T_3605; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_13 = _T_3614; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_14 = _T_3623; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_15 = _T_3632; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_16 = _T_3641; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_17 = _T_3650; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_18 = _T_3659; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_19 = _T_3668; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_20 = _T_3677; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_21 = _T_3686; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_22 = _T_3695; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_23 = _T_3704; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_24 = _T_3713; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_25 = _T_3722; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_26 = _T_3731; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_27 = _T_3740; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_28 = _T_3749; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_29 = _T_3758; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_30 = _T_3767; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_31 = _T_3776; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_32 = _T_3785; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_33 = _T_3794; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_34 = _T_3803; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_35 = _T_3812; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_36 = _T_3821; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_37 = _T_3830; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_38 = _T_3839; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_39 = _T_3848; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_40 = _T_3857; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_41 = _T_3866; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_42 = _T_3875; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_43 = _T_3884; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_44 = _T_3893; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_45 = _T_3902; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_46 = _T_3911; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_47 = _T_3920; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_48 = _T_3929; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_49 = _T_3938; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_50 = _T_3947; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_51 = _T_3956; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_52 = _T_3965; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_53 = _T_3974; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_54 = _T_3983; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_55 = _T_3992; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_56 = _T_4001; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_57 = _T_4010; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_58 = _T_4019; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_59 = _T_4028; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_60 = _T_4037; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_61 = _T_4046; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_62 = _T_4055; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_63 = _T_4064; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_64 = _T_4073; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_65 = _T_4082; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_66 = _T_4091; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_67 = _T_4100; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_68 = _T_4109; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_69 = _T_4118; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_70 = _T_4127; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_71 = _T_4136; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_72 = _T_4145; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_73 = _T_4154; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_74 = _T_4163; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_75 = _T_4172; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_76 = _T_4181; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_77 = _T_4190; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_78 = _T_4199; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_79 = _T_4208; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_80 = _T_4217; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_81 = _T_4226; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_82 = _T_4235; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_83 = _T_4244; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_84 = _T_4253; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_85 = _T_4262; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_86 = _T_4271; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_87 = _T_4280; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_88 = _T_4289; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_89 = _T_4298; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_90 = _T_4307; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_91 = _T_4316; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_92 = _T_4325; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_93 = _T_4334; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_94 = _T_4343; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_95 = _T_4352; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_96 = _T_4361; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_97 = _T_4370; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_98 = _T_4379; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_99 = _T_4388; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_100 = _T_4397; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_101 = _T_4406; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_102 = _T_4415; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_103 = _T_4424; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_104 = _T_4433; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_105 = _T_4442; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_106 = _T_4451; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_107 = _T_4460; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_108 = _T_4469; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_109 = _T_4478; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_110 = _T_4487; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_111 = _T_4496; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_112 = _T_4505; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_113 = _T_4514; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_114 = _T_4523; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_115 = _T_4532; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_116 = _T_4541; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_117 = _T_4550; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_118 = _T_4559; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_119 = _T_4568; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_120 = _T_4577; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_121 = _T_4586; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_122 = _T_4595; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_123 = _T_4604; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_124 = _T_4613; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_125 = _T_4622; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_126 = _T_4631; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_dataInput_127 = _T_4640; // @[GraphicEngineVGA.scala 308:50]
  assign multiHotPriortyReductionTree_io_selectInput_0 = _T_3500 & _T_3503; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_1 = _T_3509 & _T_3512; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_2 = _T_3518 & _T_3521; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_3 = _T_3527 & _T_3530; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_4 = _T_3536 & _T_3539; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_5 = _T_3545 & _T_3548; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_6 = _T_3554 & _T_3557; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_7 = _T_3563 & _T_3566; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_8 = _T_3572 & _T_3575; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_9 = _T_3581 & _T_3584; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_10 = _T_3590 & _T_3593; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_11 = _T_3599 & _T_3602; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_12 = _T_3608 & _T_3611; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_13 = _T_3617 & _T_3620; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_14 = _T_3626 & _T_3629; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_15 = _T_3635 & _T_3638; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_16 = _T_3644 & _T_3647; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_17 = _T_3653 & _T_3656; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_18 = _T_3662 & _T_3665; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_19 = _T_3671 & _T_3674; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_20 = _T_3680 & _T_3683; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_21 = _T_3689 & _T_3692; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_22 = _T_3698 & _T_3701; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_23 = _T_3707 & _T_3710; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_24 = _T_3716 & _T_3719; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_25 = _T_3725 & _T_3728; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_26 = _T_3734 & _T_3737; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_27 = _T_3743 & _T_3746; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_28 = _T_3752 & _T_3755; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_29 = _T_3761 & _T_3764; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_30 = _T_3770 & _T_3773; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_31 = _T_3779 & _T_3782; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_32 = _T_3788 & _T_3791; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_33 = _T_3797 & _T_3800; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_34 = _T_3805_0 & _T_3809; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_35 = _T_3814_0 & _T_3818; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_36 = _T_3823_0 & _T_3827; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_37 = _T_3832_0 & _T_3836; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_38 = _T_3841_0 & _T_3845; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_39 = _T_3850_0 & _T_3854; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_40 = _T_3859_0 & _T_3863; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_41 = _T_3869 & _T_3872; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_42 = _T_3878 & _T_3881; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_43 = _T_3887 & _T_3890; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_44 = _T_3896 & _T_3899; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_45 = _T_3905 & _T_3908; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_46 = _T_3914 & _T_3917; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_47 = _T_3923 & _T_3926; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_48 = _T_3932 & _T_3935; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_49 = _T_3941 & _T_3944; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_50 = _T_3950 & _T_3953; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_51 = _T_3959 & _T_3962; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_52 = _T_3967_0 & _T_3971; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_53 = _T_3976_0 & _T_3980; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_54 = _T_3985_0 & _T_3989; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_55 = _T_3995 & _T_3998; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_56 = _T_4004 & _T_4007; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_57 = _T_4013 & _T_4016; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_58 = _T_4021_0 & _T_4025; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_59 = _T_4030_0 & _T_4034; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_60 = _T_4039_0 & _T_4043; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_61 = _T_4049 & _T_4052; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_62 = _T_4058 & _T_4061; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_63 = _T_4067 & _T_4070; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_64 = _T_4076 & _T_4079; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_65 = _T_4085 & _T_4088; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_66 = _T_4094 & _T_4097; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_67 = _T_4102_0 & _T_4106; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_68 = _T_4111_0 & _T_4115; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_69 = _T_4120_0 & _T_4124; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_70 = _T_4130 & _T_4133; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_71 = _T_4139 & _T_4142; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_72 = _T_4148 & _T_4151; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_73 = _T_4156_0 & _T_4160; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_74 = _T_4165_0 & _T_4169; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_75 = _T_4174_0 & _T_4178; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_76 = _T_4183_0 & _T_4187; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_77 = _T_4192_0 & _T_4196; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_78 = _T_4201_0 & _T_4205; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_79 = _T_4210_0 & _T_4214; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_80 = _T_4219_0 & _T_4223; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_81 = _T_4228_0 & _T_4232; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_82 = _T_4237_0 & _T_4241; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_83 = _T_4246_0 & _T_4250; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_84 = _T_4255_0 & _T_4259; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_85 = _T_4264_0 & _T_4268; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_86 = _T_4273_0 & _T_4277; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_87 = _T_4282_0 & _T_4286; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_88 = _T_4291_0 & _T_4295; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_89 = _T_4300_0 & _T_4304; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_90 = _T_4309_0 & _T_4313; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_91 = _T_4318_0 & _T_4322; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_92 = _T_4327_0 & _T_4331; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_93 = _T_4336_0 & _T_4340; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_94 = _T_4345_0 & _T_4349; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_95 = _T_4354_0 & _T_4358; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_96 = _T_4363_0 & _T_4367; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_97 = _T_4372_0 & _T_4376; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_98 = _T_4381_0 & _T_4385; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_99 = _T_4390_0 & _T_4394; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_100 = _T_4399_0 & _T_4403; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_101 = _T_4408_0 & _T_4412; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_102 = _T_4417_0 & _T_4421; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_103 = _T_4426_0 & _T_4430; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_104 = _T_4435_0 & _T_4439; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_105 = _T_4444_0 & _T_4448; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_106 = _T_4453_0 & _T_4457; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_107 = _T_4462_0 & _T_4466; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_108 = _T_4471_0 & _T_4475; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_109 = _T_4480_0 & _T_4484; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_110 = _T_4489_0 & _T_4493; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_111 = _T_4498_0 & _T_4502; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_112 = _T_4507_0 & _T_4511; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_113 = _T_4516_0 & _T_4520; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_114 = _T_4525_0 & _T_4529; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_115 = _T_4534_0 & _T_4538; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_116 = _T_4543_0 & _T_4547; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_117 = _T_4552_0 & _T_4556; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_118 = _T_4561_0 & _T_4565; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_119 = _T_4570_0 & _T_4574; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_120 = _T_4579_0 & _T_4583; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_121 = _T_4588_0 & _T_4592; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_122 = _T_4597_0 & _T_4601; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_123 = _T_4606_0 & _T_4610; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_124 = _T_4615_0 & _T_4619; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_125 = _T_4624_0 & _T_4628; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_126 = _T_4633_0 & _T_4637; // @[GraphicEngineVGA.scala 309:52]
  assign multiHotPriortyReductionTree_io_selectInput_127 = _T_4642_0 & _T_4646; // @[GraphicEngineVGA.scala 309:52]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ScaleCounterReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  CounterXReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  CounterYReg = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  backMemoryRestoreCounter = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  _T_14_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_14_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_14_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_14_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_16_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_16_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_16_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_16_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  frameClockCount = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  spriteXPositionReg_0 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  spriteXPositionReg_1 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  spriteXPositionReg_2 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  spriteXPositionReg_3 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  spriteXPositionReg_4 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  spriteXPositionReg_5 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  spriteXPositionReg_6 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  spriteXPositionReg_7 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  spriteXPositionReg_8 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  spriteXPositionReg_9 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  spriteXPositionReg_10 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  spriteXPositionReg_11 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  spriteXPositionReg_12 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  spriteXPositionReg_13 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  spriteXPositionReg_14 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  spriteXPositionReg_15 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  spriteXPositionReg_16 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  spriteXPositionReg_17 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  spriteXPositionReg_18 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  spriteXPositionReg_19 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  spriteXPositionReg_20 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  spriteXPositionReg_21 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  spriteXPositionReg_22 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  spriteXPositionReg_23 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  spriteXPositionReg_24 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  spriteXPositionReg_25 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  spriteXPositionReg_26 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  spriteXPositionReg_27 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  spriteXPositionReg_28 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  spriteXPositionReg_29 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  spriteXPositionReg_30 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  spriteXPositionReg_31 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  spriteXPositionReg_32 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  spriteXPositionReg_33 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  spriteXPositionReg_34 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  spriteXPositionReg_35 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  spriteXPositionReg_36 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  spriteXPositionReg_37 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  spriteXPositionReg_38 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  spriteXPositionReg_39 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  spriteXPositionReg_40 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  spriteXPositionReg_41 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  spriteXPositionReg_42 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  spriteXPositionReg_43 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  spriteXPositionReg_44 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  spriteXPositionReg_45 = _RAND_58[10:0];
  _RAND_59 = {1{`RANDOM}};
  spriteXPositionReg_46 = _RAND_59[10:0];
  _RAND_60 = {1{`RANDOM}};
  spriteXPositionReg_47 = _RAND_60[10:0];
  _RAND_61 = {1{`RANDOM}};
  spriteXPositionReg_48 = _RAND_61[10:0];
  _RAND_62 = {1{`RANDOM}};
  spriteXPositionReg_49 = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  spriteXPositionReg_50 = _RAND_63[10:0];
  _RAND_64 = {1{`RANDOM}};
  spriteXPositionReg_51 = _RAND_64[10:0];
  _RAND_65 = {1{`RANDOM}};
  spriteXPositionReg_52 = _RAND_65[10:0];
  _RAND_66 = {1{`RANDOM}};
  spriteXPositionReg_53 = _RAND_66[10:0];
  _RAND_67 = {1{`RANDOM}};
  spriteXPositionReg_54 = _RAND_67[10:0];
  _RAND_68 = {1{`RANDOM}};
  spriteXPositionReg_55 = _RAND_68[10:0];
  _RAND_69 = {1{`RANDOM}};
  spriteXPositionReg_56 = _RAND_69[10:0];
  _RAND_70 = {1{`RANDOM}};
  spriteXPositionReg_57 = _RAND_70[10:0];
  _RAND_71 = {1{`RANDOM}};
  spriteXPositionReg_58 = _RAND_71[10:0];
  _RAND_72 = {1{`RANDOM}};
  spriteXPositionReg_59 = _RAND_72[10:0];
  _RAND_73 = {1{`RANDOM}};
  spriteXPositionReg_60 = _RAND_73[10:0];
  _RAND_74 = {1{`RANDOM}};
  spriteXPositionReg_61 = _RAND_74[10:0];
  _RAND_75 = {1{`RANDOM}};
  spriteXPositionReg_62 = _RAND_75[10:0];
  _RAND_76 = {1{`RANDOM}};
  spriteXPositionReg_63 = _RAND_76[10:0];
  _RAND_77 = {1{`RANDOM}};
  spriteXPositionReg_64 = _RAND_77[10:0];
  _RAND_78 = {1{`RANDOM}};
  spriteXPositionReg_65 = _RAND_78[10:0];
  _RAND_79 = {1{`RANDOM}};
  spriteXPositionReg_66 = _RAND_79[10:0];
  _RAND_80 = {1{`RANDOM}};
  spriteXPositionReg_67 = _RAND_80[10:0];
  _RAND_81 = {1{`RANDOM}};
  spriteXPositionReg_68 = _RAND_81[10:0];
  _RAND_82 = {1{`RANDOM}};
  spriteXPositionReg_69 = _RAND_82[10:0];
  _RAND_83 = {1{`RANDOM}};
  spriteXPositionReg_70 = _RAND_83[10:0];
  _RAND_84 = {1{`RANDOM}};
  spriteXPositionReg_71 = _RAND_84[10:0];
  _RAND_85 = {1{`RANDOM}};
  spriteXPositionReg_72 = _RAND_85[10:0];
  _RAND_86 = {1{`RANDOM}};
  spriteXPositionReg_73 = _RAND_86[10:0];
  _RAND_87 = {1{`RANDOM}};
  spriteXPositionReg_74 = _RAND_87[10:0];
  _RAND_88 = {1{`RANDOM}};
  spriteXPositionReg_75 = _RAND_88[10:0];
  _RAND_89 = {1{`RANDOM}};
  spriteXPositionReg_76 = _RAND_89[10:0];
  _RAND_90 = {1{`RANDOM}};
  spriteXPositionReg_77 = _RAND_90[10:0];
  _RAND_91 = {1{`RANDOM}};
  spriteXPositionReg_78 = _RAND_91[10:0];
  _RAND_92 = {1{`RANDOM}};
  spriteXPositionReg_79 = _RAND_92[10:0];
  _RAND_93 = {1{`RANDOM}};
  spriteXPositionReg_80 = _RAND_93[10:0];
  _RAND_94 = {1{`RANDOM}};
  spriteXPositionReg_81 = _RAND_94[10:0];
  _RAND_95 = {1{`RANDOM}};
  spriteXPositionReg_82 = _RAND_95[10:0];
  _RAND_96 = {1{`RANDOM}};
  spriteXPositionReg_83 = _RAND_96[10:0];
  _RAND_97 = {1{`RANDOM}};
  spriteXPositionReg_84 = _RAND_97[10:0];
  _RAND_98 = {1{`RANDOM}};
  spriteXPositionReg_85 = _RAND_98[10:0];
  _RAND_99 = {1{`RANDOM}};
  spriteXPositionReg_86 = _RAND_99[10:0];
  _RAND_100 = {1{`RANDOM}};
  spriteXPositionReg_87 = _RAND_100[10:0];
  _RAND_101 = {1{`RANDOM}};
  spriteXPositionReg_88 = _RAND_101[10:0];
  _RAND_102 = {1{`RANDOM}};
  spriteXPositionReg_89 = _RAND_102[10:0];
  _RAND_103 = {1{`RANDOM}};
  spriteXPositionReg_90 = _RAND_103[10:0];
  _RAND_104 = {1{`RANDOM}};
  spriteXPositionReg_91 = _RAND_104[10:0];
  _RAND_105 = {1{`RANDOM}};
  spriteXPositionReg_92 = _RAND_105[10:0];
  _RAND_106 = {1{`RANDOM}};
  spriteXPositionReg_93 = _RAND_106[10:0];
  _RAND_107 = {1{`RANDOM}};
  spriteXPositionReg_94 = _RAND_107[10:0];
  _RAND_108 = {1{`RANDOM}};
  spriteXPositionReg_95 = _RAND_108[10:0];
  _RAND_109 = {1{`RANDOM}};
  spriteXPositionReg_96 = _RAND_109[10:0];
  _RAND_110 = {1{`RANDOM}};
  spriteXPositionReg_97 = _RAND_110[10:0];
  _RAND_111 = {1{`RANDOM}};
  spriteXPositionReg_98 = _RAND_111[10:0];
  _RAND_112 = {1{`RANDOM}};
  spriteXPositionReg_99 = _RAND_112[10:0];
  _RAND_113 = {1{`RANDOM}};
  spriteXPositionReg_100 = _RAND_113[10:0];
  _RAND_114 = {1{`RANDOM}};
  spriteXPositionReg_101 = _RAND_114[10:0];
  _RAND_115 = {1{`RANDOM}};
  spriteXPositionReg_102 = _RAND_115[10:0];
  _RAND_116 = {1{`RANDOM}};
  spriteXPositionReg_103 = _RAND_116[10:0];
  _RAND_117 = {1{`RANDOM}};
  spriteXPositionReg_104 = _RAND_117[10:0];
  _RAND_118 = {1{`RANDOM}};
  spriteXPositionReg_105 = _RAND_118[10:0];
  _RAND_119 = {1{`RANDOM}};
  spriteXPositionReg_106 = _RAND_119[10:0];
  _RAND_120 = {1{`RANDOM}};
  spriteXPositionReg_107 = _RAND_120[10:0];
  _RAND_121 = {1{`RANDOM}};
  spriteXPositionReg_108 = _RAND_121[10:0];
  _RAND_122 = {1{`RANDOM}};
  spriteXPositionReg_109 = _RAND_122[10:0];
  _RAND_123 = {1{`RANDOM}};
  spriteXPositionReg_110 = _RAND_123[10:0];
  _RAND_124 = {1{`RANDOM}};
  spriteXPositionReg_111 = _RAND_124[10:0];
  _RAND_125 = {1{`RANDOM}};
  spriteXPositionReg_112 = _RAND_125[10:0];
  _RAND_126 = {1{`RANDOM}};
  spriteXPositionReg_113 = _RAND_126[10:0];
  _RAND_127 = {1{`RANDOM}};
  spriteXPositionReg_114 = _RAND_127[10:0];
  _RAND_128 = {1{`RANDOM}};
  spriteXPositionReg_115 = _RAND_128[10:0];
  _RAND_129 = {1{`RANDOM}};
  spriteXPositionReg_116 = _RAND_129[10:0];
  _RAND_130 = {1{`RANDOM}};
  spriteXPositionReg_117 = _RAND_130[10:0];
  _RAND_131 = {1{`RANDOM}};
  spriteXPositionReg_118 = _RAND_131[10:0];
  _RAND_132 = {1{`RANDOM}};
  spriteXPositionReg_119 = _RAND_132[10:0];
  _RAND_133 = {1{`RANDOM}};
  spriteXPositionReg_120 = _RAND_133[10:0];
  _RAND_134 = {1{`RANDOM}};
  spriteXPositionReg_121 = _RAND_134[10:0];
  _RAND_135 = {1{`RANDOM}};
  spriteXPositionReg_122 = _RAND_135[10:0];
  _RAND_136 = {1{`RANDOM}};
  spriteXPositionReg_123 = _RAND_136[10:0];
  _RAND_137 = {1{`RANDOM}};
  spriteXPositionReg_124 = _RAND_137[10:0];
  _RAND_138 = {1{`RANDOM}};
  spriteXPositionReg_125 = _RAND_138[10:0];
  _RAND_139 = {1{`RANDOM}};
  spriteXPositionReg_126 = _RAND_139[10:0];
  _RAND_140 = {1{`RANDOM}};
  spriteXPositionReg_127 = _RAND_140[10:0];
  _RAND_141 = {1{`RANDOM}};
  spriteYPositionReg_0 = _RAND_141[9:0];
  _RAND_142 = {1{`RANDOM}};
  spriteYPositionReg_1 = _RAND_142[9:0];
  _RAND_143 = {1{`RANDOM}};
  spriteYPositionReg_2 = _RAND_143[9:0];
  _RAND_144 = {1{`RANDOM}};
  spriteYPositionReg_3 = _RAND_144[9:0];
  _RAND_145 = {1{`RANDOM}};
  spriteYPositionReg_4 = _RAND_145[9:0];
  _RAND_146 = {1{`RANDOM}};
  spriteYPositionReg_5 = _RAND_146[9:0];
  _RAND_147 = {1{`RANDOM}};
  spriteYPositionReg_6 = _RAND_147[9:0];
  _RAND_148 = {1{`RANDOM}};
  spriteYPositionReg_7 = _RAND_148[9:0];
  _RAND_149 = {1{`RANDOM}};
  spriteYPositionReg_8 = _RAND_149[9:0];
  _RAND_150 = {1{`RANDOM}};
  spriteYPositionReg_9 = _RAND_150[9:0];
  _RAND_151 = {1{`RANDOM}};
  spriteYPositionReg_10 = _RAND_151[9:0];
  _RAND_152 = {1{`RANDOM}};
  spriteYPositionReg_11 = _RAND_152[9:0];
  _RAND_153 = {1{`RANDOM}};
  spriteYPositionReg_12 = _RAND_153[9:0];
  _RAND_154 = {1{`RANDOM}};
  spriteYPositionReg_13 = _RAND_154[9:0];
  _RAND_155 = {1{`RANDOM}};
  spriteYPositionReg_14 = _RAND_155[9:0];
  _RAND_156 = {1{`RANDOM}};
  spriteYPositionReg_15 = _RAND_156[9:0];
  _RAND_157 = {1{`RANDOM}};
  spriteYPositionReg_16 = _RAND_157[9:0];
  _RAND_158 = {1{`RANDOM}};
  spriteYPositionReg_17 = _RAND_158[9:0];
  _RAND_159 = {1{`RANDOM}};
  spriteYPositionReg_18 = _RAND_159[9:0];
  _RAND_160 = {1{`RANDOM}};
  spriteYPositionReg_19 = _RAND_160[9:0];
  _RAND_161 = {1{`RANDOM}};
  spriteYPositionReg_20 = _RAND_161[9:0];
  _RAND_162 = {1{`RANDOM}};
  spriteYPositionReg_21 = _RAND_162[9:0];
  _RAND_163 = {1{`RANDOM}};
  spriteYPositionReg_22 = _RAND_163[9:0];
  _RAND_164 = {1{`RANDOM}};
  spriteYPositionReg_23 = _RAND_164[9:0];
  _RAND_165 = {1{`RANDOM}};
  spriteYPositionReg_24 = _RAND_165[9:0];
  _RAND_166 = {1{`RANDOM}};
  spriteYPositionReg_25 = _RAND_166[9:0];
  _RAND_167 = {1{`RANDOM}};
  spriteYPositionReg_26 = _RAND_167[9:0];
  _RAND_168 = {1{`RANDOM}};
  spriteYPositionReg_27 = _RAND_168[9:0];
  _RAND_169 = {1{`RANDOM}};
  spriteYPositionReg_28 = _RAND_169[9:0];
  _RAND_170 = {1{`RANDOM}};
  spriteYPositionReg_29 = _RAND_170[9:0];
  _RAND_171 = {1{`RANDOM}};
  spriteYPositionReg_30 = _RAND_171[9:0];
  _RAND_172 = {1{`RANDOM}};
  spriteYPositionReg_31 = _RAND_172[9:0];
  _RAND_173 = {1{`RANDOM}};
  spriteYPositionReg_32 = _RAND_173[9:0];
  _RAND_174 = {1{`RANDOM}};
  spriteYPositionReg_33 = _RAND_174[9:0];
  _RAND_175 = {1{`RANDOM}};
  spriteYPositionReg_34 = _RAND_175[9:0];
  _RAND_176 = {1{`RANDOM}};
  spriteYPositionReg_35 = _RAND_176[9:0];
  _RAND_177 = {1{`RANDOM}};
  spriteYPositionReg_36 = _RAND_177[9:0];
  _RAND_178 = {1{`RANDOM}};
  spriteYPositionReg_37 = _RAND_178[9:0];
  _RAND_179 = {1{`RANDOM}};
  spriteYPositionReg_38 = _RAND_179[9:0];
  _RAND_180 = {1{`RANDOM}};
  spriteYPositionReg_39 = _RAND_180[9:0];
  _RAND_181 = {1{`RANDOM}};
  spriteYPositionReg_40 = _RAND_181[9:0];
  _RAND_182 = {1{`RANDOM}};
  spriteYPositionReg_41 = _RAND_182[9:0];
  _RAND_183 = {1{`RANDOM}};
  spriteYPositionReg_42 = _RAND_183[9:0];
  _RAND_184 = {1{`RANDOM}};
  spriteYPositionReg_43 = _RAND_184[9:0];
  _RAND_185 = {1{`RANDOM}};
  spriteYPositionReg_44 = _RAND_185[9:0];
  _RAND_186 = {1{`RANDOM}};
  spriteYPositionReg_45 = _RAND_186[9:0];
  _RAND_187 = {1{`RANDOM}};
  spriteYPositionReg_46 = _RAND_187[9:0];
  _RAND_188 = {1{`RANDOM}};
  spriteYPositionReg_47 = _RAND_188[9:0];
  _RAND_189 = {1{`RANDOM}};
  spriteYPositionReg_48 = _RAND_189[9:0];
  _RAND_190 = {1{`RANDOM}};
  spriteYPositionReg_49 = _RAND_190[9:0];
  _RAND_191 = {1{`RANDOM}};
  spriteYPositionReg_50 = _RAND_191[9:0];
  _RAND_192 = {1{`RANDOM}};
  spriteYPositionReg_51 = _RAND_192[9:0];
  _RAND_193 = {1{`RANDOM}};
  spriteYPositionReg_52 = _RAND_193[9:0];
  _RAND_194 = {1{`RANDOM}};
  spriteYPositionReg_53 = _RAND_194[9:0];
  _RAND_195 = {1{`RANDOM}};
  spriteYPositionReg_54 = _RAND_195[9:0];
  _RAND_196 = {1{`RANDOM}};
  spriteYPositionReg_55 = _RAND_196[9:0];
  _RAND_197 = {1{`RANDOM}};
  spriteYPositionReg_56 = _RAND_197[9:0];
  _RAND_198 = {1{`RANDOM}};
  spriteYPositionReg_57 = _RAND_198[9:0];
  _RAND_199 = {1{`RANDOM}};
  spriteYPositionReg_58 = _RAND_199[9:0];
  _RAND_200 = {1{`RANDOM}};
  spriteYPositionReg_59 = _RAND_200[9:0];
  _RAND_201 = {1{`RANDOM}};
  spriteYPositionReg_60 = _RAND_201[9:0];
  _RAND_202 = {1{`RANDOM}};
  spriteYPositionReg_61 = _RAND_202[9:0];
  _RAND_203 = {1{`RANDOM}};
  spriteYPositionReg_62 = _RAND_203[9:0];
  _RAND_204 = {1{`RANDOM}};
  spriteYPositionReg_63 = _RAND_204[9:0];
  _RAND_205 = {1{`RANDOM}};
  spriteYPositionReg_70 = _RAND_205[9:0];
  _RAND_206 = {1{`RANDOM}};
  spriteYPositionReg_71 = _RAND_206[9:0];
  _RAND_207 = {1{`RANDOM}};
  spriteYPositionReg_72 = _RAND_207[9:0];
  _RAND_208 = {1{`RANDOM}};
  spriteYPositionReg_73 = _RAND_208[9:0];
  _RAND_209 = {1{`RANDOM}};
  spriteYPositionReg_74 = _RAND_209[9:0];
  _RAND_210 = {1{`RANDOM}};
  spriteYPositionReg_75 = _RAND_210[9:0];
  _RAND_211 = {1{`RANDOM}};
  spriteYPositionReg_76 = _RAND_211[9:0];
  _RAND_212 = {1{`RANDOM}};
  spriteYPositionReg_77 = _RAND_212[9:0];
  _RAND_213 = {1{`RANDOM}};
  spriteYPositionReg_78 = _RAND_213[9:0];
  _RAND_214 = {1{`RANDOM}};
  spriteYPositionReg_79 = _RAND_214[9:0];
  _RAND_215 = {1{`RANDOM}};
  spriteYPositionReg_80 = _RAND_215[9:0];
  _RAND_216 = {1{`RANDOM}};
  spriteYPositionReg_81 = _RAND_216[9:0];
  _RAND_217 = {1{`RANDOM}};
  spriteYPositionReg_82 = _RAND_217[9:0];
  _RAND_218 = {1{`RANDOM}};
  spriteYPositionReg_83 = _RAND_218[9:0];
  _RAND_219 = {1{`RANDOM}};
  spriteYPositionReg_84 = _RAND_219[9:0];
  _RAND_220 = {1{`RANDOM}};
  spriteYPositionReg_85 = _RAND_220[9:0];
  _RAND_221 = {1{`RANDOM}};
  spriteYPositionReg_86 = _RAND_221[9:0];
  _RAND_222 = {1{`RANDOM}};
  spriteYPositionReg_87 = _RAND_222[9:0];
  _RAND_223 = {1{`RANDOM}};
  spriteYPositionReg_88 = _RAND_223[9:0];
  _RAND_224 = {1{`RANDOM}};
  spriteYPositionReg_89 = _RAND_224[9:0];
  _RAND_225 = {1{`RANDOM}};
  spriteYPositionReg_90 = _RAND_225[9:0];
  _RAND_226 = {1{`RANDOM}};
  spriteYPositionReg_91 = _RAND_226[9:0];
  _RAND_227 = {1{`RANDOM}};
  spriteYPositionReg_92 = _RAND_227[9:0];
  _RAND_228 = {1{`RANDOM}};
  spriteYPositionReg_93 = _RAND_228[9:0];
  _RAND_229 = {1{`RANDOM}};
  spriteYPositionReg_94 = _RAND_229[9:0];
  _RAND_230 = {1{`RANDOM}};
  spriteYPositionReg_95 = _RAND_230[9:0];
  _RAND_231 = {1{`RANDOM}};
  spriteYPositionReg_96 = _RAND_231[9:0];
  _RAND_232 = {1{`RANDOM}};
  spriteYPositionReg_97 = _RAND_232[9:0];
  _RAND_233 = {1{`RANDOM}};
  spriteYPositionReg_98 = _RAND_233[9:0];
  _RAND_234 = {1{`RANDOM}};
  spriteYPositionReg_99 = _RAND_234[9:0];
  _RAND_235 = {1{`RANDOM}};
  spriteYPositionReg_100 = _RAND_235[9:0];
  _RAND_236 = {1{`RANDOM}};
  spriteYPositionReg_101 = _RAND_236[9:0];
  _RAND_237 = {1{`RANDOM}};
  spriteYPositionReg_102 = _RAND_237[9:0];
  _RAND_238 = {1{`RANDOM}};
  spriteYPositionReg_103 = _RAND_238[9:0];
  _RAND_239 = {1{`RANDOM}};
  spriteYPositionReg_104 = _RAND_239[9:0];
  _RAND_240 = {1{`RANDOM}};
  spriteYPositionReg_105 = _RAND_240[9:0];
  _RAND_241 = {1{`RANDOM}};
  spriteYPositionReg_106 = _RAND_241[9:0];
  _RAND_242 = {1{`RANDOM}};
  spriteYPositionReg_107 = _RAND_242[9:0];
  _RAND_243 = {1{`RANDOM}};
  spriteYPositionReg_108 = _RAND_243[9:0];
  _RAND_244 = {1{`RANDOM}};
  spriteYPositionReg_109 = _RAND_244[9:0];
  _RAND_245 = {1{`RANDOM}};
  spriteYPositionReg_110 = _RAND_245[9:0];
  _RAND_246 = {1{`RANDOM}};
  spriteYPositionReg_111 = _RAND_246[9:0];
  _RAND_247 = {1{`RANDOM}};
  spriteYPositionReg_112 = _RAND_247[9:0];
  _RAND_248 = {1{`RANDOM}};
  spriteYPositionReg_113 = _RAND_248[9:0];
  _RAND_249 = {1{`RANDOM}};
  spriteYPositionReg_114 = _RAND_249[9:0];
  _RAND_250 = {1{`RANDOM}};
  spriteYPositionReg_115 = _RAND_250[9:0];
  _RAND_251 = {1{`RANDOM}};
  spriteYPositionReg_116 = _RAND_251[9:0];
  _RAND_252 = {1{`RANDOM}};
  spriteYPositionReg_117 = _RAND_252[9:0];
  _RAND_253 = {1{`RANDOM}};
  spriteYPositionReg_118 = _RAND_253[9:0];
  _RAND_254 = {1{`RANDOM}};
  spriteYPositionReg_119 = _RAND_254[9:0];
  _RAND_255 = {1{`RANDOM}};
  spriteYPositionReg_120 = _RAND_255[9:0];
  _RAND_256 = {1{`RANDOM}};
  spriteYPositionReg_121 = _RAND_256[9:0];
  _RAND_257 = {1{`RANDOM}};
  spriteYPositionReg_122 = _RAND_257[9:0];
  _RAND_258 = {1{`RANDOM}};
  spriteYPositionReg_123 = _RAND_258[9:0];
  _RAND_259 = {1{`RANDOM}};
  spriteYPositionReg_124 = _RAND_259[9:0];
  _RAND_260 = {1{`RANDOM}};
  spriteYPositionReg_125 = _RAND_260[9:0];
  _RAND_261 = {1{`RANDOM}};
  spriteYPositionReg_126 = _RAND_261[9:0];
  _RAND_262 = {1{`RANDOM}};
  spriteYPositionReg_127 = _RAND_262[9:0];
  _RAND_263 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  spriteVisibleReg_32 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  spriteVisibleReg_33 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  spriteVisibleReg_41 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  spriteVisibleReg_42 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  spriteVisibleReg_43 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  spriteVisibleReg_44 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  spriteVisibleReg_45 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  spriteVisibleReg_46 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  spriteVisibleReg_47 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  spriteVisibleReg_48 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  spriteVisibleReg_49 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  spriteVisibleReg_50 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  spriteVisibleReg_51 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  spriteVisibleReg_55 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  spriteVisibleReg_56 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  spriteVisibleReg_57 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  spriteVisibleReg_61 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  spriteVisibleReg_62 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  spriteVisibleReg_63 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  spriteVisibleReg_64 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  spriteVisibleReg_65 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  spriteVisibleReg_66 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  spriteVisibleReg_70 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  spriteVisibleReg_71 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  spriteVisibleReg_72 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  spriteFlipVerticalReg_122 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  spriteFlipVerticalReg_123 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  spriteFlipVerticalReg_124 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  spriteFlipVerticalReg_125 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  spriteFlipVerticalReg_126 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  spriteFlipVerticalReg_127 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  viewBoxXReg_0 = _RAND_326[9:0];
  _RAND_327 = {1{`RANDOM}};
  missingFrameErrorReg = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  backBufferWriteErrorReg = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  viewBoxOutOfRangeErrorReg = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  newFrameStikyReg = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  _T_43 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  backTileMemoryDataRead_0_0 = _RAND_332[6:0];
  _RAND_333 = {1{`RANDOM}};
  backTileMemoryDataRead_0_1 = _RAND_333[6:0];
  _RAND_334 = {1{`RANDOM}};
  backTileMemoryDataRead_0_2 = _RAND_334[6:0];
  _RAND_335 = {1{`RANDOM}};
  backTileMemoryDataRead_0_3 = _RAND_335[6:0];
  _RAND_336 = {1{`RANDOM}};
  backTileMemoryDataRead_0_4 = _RAND_336[6:0];
  _RAND_337 = {1{`RANDOM}};
  backTileMemoryDataRead_0_5 = _RAND_337[6:0];
  _RAND_338 = {1{`RANDOM}};
  backTileMemoryDataRead_0_6 = _RAND_338[6:0];
  _RAND_339 = {1{`RANDOM}};
  backTileMemoryDataRead_0_7 = _RAND_339[6:0];
  _RAND_340 = {1{`RANDOM}};
  backTileMemoryDataRead_0_8 = _RAND_340[6:0];
  _RAND_341 = {1{`RANDOM}};
  backTileMemoryDataRead_0_9 = _RAND_341[6:0];
  _RAND_342 = {1{`RANDOM}};
  backTileMemoryDataRead_0_10 = _RAND_342[6:0];
  _RAND_343 = {1{`RANDOM}};
  backTileMemoryDataRead_0_11 = _RAND_343[6:0];
  _RAND_344 = {1{`RANDOM}};
  backTileMemoryDataRead_0_12 = _RAND_344[6:0];
  _RAND_345 = {1{`RANDOM}};
  backTileMemoryDataRead_0_13 = _RAND_345[6:0];
  _RAND_346 = {1{`RANDOM}};
  backTileMemoryDataRead_0_14 = _RAND_346[6:0];
  _RAND_347 = {1{`RANDOM}};
  backTileMemoryDataRead_0_15 = _RAND_347[6:0];
  _RAND_348 = {1{`RANDOM}};
  backTileMemoryDataRead_0_16 = _RAND_348[6:0];
  _RAND_349 = {1{`RANDOM}};
  backTileMemoryDataRead_0_17 = _RAND_349[6:0];
  _RAND_350 = {1{`RANDOM}};
  backTileMemoryDataRead_0_18 = _RAND_350[6:0];
  _RAND_351 = {1{`RANDOM}};
  backTileMemoryDataRead_0_19 = _RAND_351[6:0];
  _RAND_352 = {1{`RANDOM}};
  backTileMemoryDataRead_0_20 = _RAND_352[6:0];
  _RAND_353 = {1{`RANDOM}};
  backTileMemoryDataRead_0_21 = _RAND_353[6:0];
  _RAND_354 = {1{`RANDOM}};
  backTileMemoryDataRead_0_22 = _RAND_354[6:0];
  _RAND_355 = {1{`RANDOM}};
  backTileMemoryDataRead_0_23 = _RAND_355[6:0];
  _RAND_356 = {1{`RANDOM}};
  backTileMemoryDataRead_0_24 = _RAND_356[6:0];
  _RAND_357 = {1{`RANDOM}};
  backTileMemoryDataRead_0_25 = _RAND_357[6:0];
  _RAND_358 = {1{`RANDOM}};
  backTileMemoryDataRead_0_26 = _RAND_358[6:0];
  _RAND_359 = {1{`RANDOM}};
  backTileMemoryDataRead_0_27 = _RAND_359[6:0];
  _RAND_360 = {1{`RANDOM}};
  backTileMemoryDataRead_0_28 = _RAND_360[6:0];
  _RAND_361 = {1{`RANDOM}};
  backTileMemoryDataRead_0_29 = _RAND_361[6:0];
  _RAND_362 = {1{`RANDOM}};
  backTileMemoryDataRead_0_30 = _RAND_362[6:0];
  _RAND_363 = {1{`RANDOM}};
  backTileMemoryDataRead_0_31 = _RAND_363[6:0];
  _RAND_364 = {1{`RANDOM}};
  backTileMemoryDataRead_1_0 = _RAND_364[6:0];
  _RAND_365 = {1{`RANDOM}};
  backTileMemoryDataRead_1_1 = _RAND_365[6:0];
  _RAND_366 = {1{`RANDOM}};
  backTileMemoryDataRead_1_2 = _RAND_366[6:0];
  _RAND_367 = {1{`RANDOM}};
  backTileMemoryDataRead_1_3 = _RAND_367[6:0];
  _RAND_368 = {1{`RANDOM}};
  backTileMemoryDataRead_1_4 = _RAND_368[6:0];
  _RAND_369 = {1{`RANDOM}};
  backTileMemoryDataRead_1_5 = _RAND_369[6:0];
  _RAND_370 = {1{`RANDOM}};
  backTileMemoryDataRead_1_6 = _RAND_370[6:0];
  _RAND_371 = {1{`RANDOM}};
  backTileMemoryDataRead_1_7 = _RAND_371[6:0];
  _RAND_372 = {1{`RANDOM}};
  backTileMemoryDataRead_1_8 = _RAND_372[6:0];
  _RAND_373 = {1{`RANDOM}};
  backTileMemoryDataRead_1_9 = _RAND_373[6:0];
  _RAND_374 = {1{`RANDOM}};
  backTileMemoryDataRead_1_10 = _RAND_374[6:0];
  _RAND_375 = {1{`RANDOM}};
  backTileMemoryDataRead_1_11 = _RAND_375[6:0];
  _RAND_376 = {1{`RANDOM}};
  backTileMemoryDataRead_1_12 = _RAND_376[6:0];
  _RAND_377 = {1{`RANDOM}};
  backTileMemoryDataRead_1_13 = _RAND_377[6:0];
  _RAND_378 = {1{`RANDOM}};
  backTileMemoryDataRead_1_14 = _RAND_378[6:0];
  _RAND_379 = {1{`RANDOM}};
  backTileMemoryDataRead_1_15 = _RAND_379[6:0];
  _RAND_380 = {1{`RANDOM}};
  backTileMemoryDataRead_1_16 = _RAND_380[6:0];
  _RAND_381 = {1{`RANDOM}};
  backTileMemoryDataRead_1_17 = _RAND_381[6:0];
  _RAND_382 = {1{`RANDOM}};
  backTileMemoryDataRead_1_18 = _RAND_382[6:0];
  _RAND_383 = {1{`RANDOM}};
  backTileMemoryDataRead_1_19 = _RAND_383[6:0];
  _RAND_384 = {1{`RANDOM}};
  backTileMemoryDataRead_1_20 = _RAND_384[6:0];
  _RAND_385 = {1{`RANDOM}};
  backTileMemoryDataRead_1_21 = _RAND_385[6:0];
  _RAND_386 = {1{`RANDOM}};
  backTileMemoryDataRead_1_22 = _RAND_386[6:0];
  _RAND_387 = {1{`RANDOM}};
  backTileMemoryDataRead_1_23 = _RAND_387[6:0];
  _RAND_388 = {1{`RANDOM}};
  backTileMemoryDataRead_1_24 = _RAND_388[6:0];
  _RAND_389 = {1{`RANDOM}};
  backTileMemoryDataRead_1_25 = _RAND_389[6:0];
  _RAND_390 = {1{`RANDOM}};
  backTileMemoryDataRead_1_26 = _RAND_390[6:0];
  _RAND_391 = {1{`RANDOM}};
  backTileMemoryDataRead_1_27 = _RAND_391[6:0];
  _RAND_392 = {1{`RANDOM}};
  backTileMemoryDataRead_1_28 = _RAND_392[6:0];
  _RAND_393 = {1{`RANDOM}};
  backTileMemoryDataRead_1_29 = _RAND_393[6:0];
  _RAND_394 = {1{`RANDOM}};
  backTileMemoryDataRead_1_30 = _RAND_394[6:0];
  _RAND_395 = {1{`RANDOM}};
  backTileMemoryDataRead_1_31 = _RAND_395[6:0];
  _RAND_396 = {1{`RANDOM}};
  backMemoryCopyCounter = _RAND_396[11:0];
  _RAND_397 = {1{`RANDOM}};
  copyEnabledReg = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  _T_373 = _RAND_398[10:0];
  _RAND_399 = {1{`RANDOM}};
  _T_375 = _RAND_399[10:0];
  _RAND_400 = {1{`RANDOM}};
  _T_378 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  _T_379 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  _T_382 = _RAND_402[4:0];
  _RAND_403 = {1{`RANDOM}};
  _T_385 = _RAND_403[10:0];
  _RAND_404 = {1{`RANDOM}};
  _T_393 = _RAND_404[10:0];
  _RAND_405 = {1{`RANDOM}};
  _T_395 = _RAND_405[10:0];
  _RAND_406 = {1{`RANDOM}};
  _T_398 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  _T_399 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  _T_402 = _RAND_408[4:0];
  _RAND_409 = {1{`RANDOM}};
  _T_405 = _RAND_409[10:0];
  _RAND_410 = {1{`RANDOM}};
  _T_412 = _RAND_410[4:0];
  _RAND_411 = {1{`RANDOM}};
  _T_415 = _RAND_411[4:0];
  _RAND_412 = {1{`RANDOM}};
  pixelColorBack = _RAND_412[5:0];
  _RAND_413 = {1{`RANDOM}};
  _T_3497 = _RAND_413[5:0];
  _RAND_414 = {1{`RANDOM}};
  _T_3498_0 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  _T_3498_1 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  _T_3499_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  _T_3499_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  _T_3502 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  _T_3506 = _RAND_419[5:0];
  _RAND_420 = {1{`RANDOM}};
  _T_3507_0 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  _T_3507_1 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  _T_3508_0 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  _T_3508_1 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  _T_3511 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  _T_3515 = _RAND_425[5:0];
  _RAND_426 = {1{`RANDOM}};
  _T_3516_0 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  _T_3516_1 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  _T_3517_0 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  _T_3517_1 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  _T_3520 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  _T_3524 = _RAND_431[5:0];
  _RAND_432 = {1{`RANDOM}};
  _T_3525_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  _T_3525_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  _T_3526_0 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  _T_3526_1 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  _T_3529 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  _T_3533 = _RAND_437[5:0];
  _RAND_438 = {1{`RANDOM}};
  _T_3534_0 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  _T_3534_1 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  _T_3535_0 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  _T_3535_1 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  _T_3538 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  _T_3542 = _RAND_443[5:0];
  _RAND_444 = {1{`RANDOM}};
  _T_3543_0 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  _T_3543_1 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  _T_3544_0 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  _T_3544_1 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  _T_3547 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  _T_3551 = _RAND_449[5:0];
  _RAND_450 = {1{`RANDOM}};
  _T_3552_0 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  _T_3552_1 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  _T_3553_0 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  _T_3553_1 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  _T_3556 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  _T_3560 = _RAND_455[5:0];
  _RAND_456 = {1{`RANDOM}};
  _T_3561_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  _T_3561_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  _T_3562_0 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  _T_3562_1 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  _T_3565 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  _T_3569 = _RAND_461[5:0];
  _RAND_462 = {1{`RANDOM}};
  _T_3570_0 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_3570_1 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_3571_0 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_3571_1 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_3574 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_3578 = _RAND_467[5:0];
  _RAND_468 = {1{`RANDOM}};
  _T_3579_0 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_3579_1 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_3580_0 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_3580_1 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_3583 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  _T_3587 = _RAND_473[5:0];
  _RAND_474 = {1{`RANDOM}};
  _T_3588_0 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  _T_3588_1 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  _T_3589_0 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  _T_3589_1 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  _T_3592 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  _T_3596 = _RAND_479[5:0];
  _RAND_480 = {1{`RANDOM}};
  _T_3597_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  _T_3597_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  _T_3598_0 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  _T_3598_1 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  _T_3601 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  _T_3605 = _RAND_485[5:0];
  _RAND_486 = {1{`RANDOM}};
  _T_3606_0 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  _T_3606_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  _T_3607_0 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  _T_3607_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  _T_3610 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  _T_3614 = _RAND_491[5:0];
  _RAND_492 = {1{`RANDOM}};
  _T_3615_0 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  _T_3615_1 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  _T_3616_0 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  _T_3616_1 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  _T_3619 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  _T_3623 = _RAND_497[5:0];
  _RAND_498 = {1{`RANDOM}};
  _T_3624_0 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  _T_3624_1 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  _T_3625_0 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  _T_3625_1 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  _T_3628 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  _T_3632 = _RAND_503[5:0];
  _RAND_504 = {1{`RANDOM}};
  _T_3633_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  _T_3633_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  _T_3634_0 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  _T_3634_1 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  _T_3637 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  _T_3641 = _RAND_509[5:0];
  _RAND_510 = {1{`RANDOM}};
  _T_3642_0 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  _T_3642_1 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  _T_3643_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  _T_3643_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  _T_3646 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  _T_3650 = _RAND_515[5:0];
  _RAND_516 = {1{`RANDOM}};
  _T_3651_0 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  _T_3651_1 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  _T_3652_0 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  _T_3652_1 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  _T_3655 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  _T_3659 = _RAND_521[5:0];
  _RAND_522 = {1{`RANDOM}};
  _T_3660_0 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  _T_3660_1 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  _T_3661_0 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  _T_3661_1 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  _T_3664 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  _T_3668 = _RAND_527[5:0];
  _RAND_528 = {1{`RANDOM}};
  _T_3669_0 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  _T_3669_1 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  _T_3670_0 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  _T_3670_1 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  _T_3673 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  _T_3677 = _RAND_533[5:0];
  _RAND_534 = {1{`RANDOM}};
  _T_3678_0 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  _T_3678_1 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  _T_3679_0 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  _T_3679_1 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  _T_3682 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  _T_3686 = _RAND_539[5:0];
  _RAND_540 = {1{`RANDOM}};
  _T_3687_0 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  _T_3687_1 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  _T_3688_0 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  _T_3688_1 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  _T_3691 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  _T_3695 = _RAND_545[5:0];
  _RAND_546 = {1{`RANDOM}};
  _T_3696_0 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  _T_3696_1 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  _T_3697_0 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  _T_3697_1 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  _T_3700 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  _T_3704 = _RAND_551[5:0];
  _RAND_552 = {1{`RANDOM}};
  _T_3705_0 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  _T_3705_1 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  _T_3706_0 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  _T_3706_1 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  _T_3709 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  _T_3713 = _RAND_557[5:0];
  _RAND_558 = {1{`RANDOM}};
  _T_3714_0 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  _T_3714_1 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  _T_3715_0 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  _T_3715_1 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  _T_3718 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  _T_3722 = _RAND_563[5:0];
  _RAND_564 = {1{`RANDOM}};
  _T_3723_0 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  _T_3723_1 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  _T_3724_0 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  _T_3724_1 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  _T_3727 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  _T_3731 = _RAND_569[5:0];
  _RAND_570 = {1{`RANDOM}};
  _T_3732_0 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  _T_3732_1 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  _T_3733_0 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  _T_3733_1 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  _T_3736 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  _T_3740 = _RAND_575[5:0];
  _RAND_576 = {1{`RANDOM}};
  _T_3741_0 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  _T_3741_1 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  _T_3742_0 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  _T_3742_1 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  _T_3745 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  _T_3749 = _RAND_581[5:0];
  _RAND_582 = {1{`RANDOM}};
  _T_3750_0 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  _T_3750_1 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  _T_3751_0 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  _T_3751_1 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  _T_3754 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  _T_3758 = _RAND_587[5:0];
  _RAND_588 = {1{`RANDOM}};
  _T_3759_0 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  _T_3759_1 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  _T_3760_0 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  _T_3760_1 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  _T_3763 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  _T_3767 = _RAND_593[5:0];
  _RAND_594 = {1{`RANDOM}};
  _T_3768_0 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  _T_3768_1 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  _T_3769_0 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  _T_3769_1 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  _T_3772 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  _T_3776 = _RAND_599[5:0];
  _RAND_600 = {1{`RANDOM}};
  _T_3777_0 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  _T_3777_1 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  _T_3778_0 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  _T_3778_1 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  _T_3781 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  _T_3785 = _RAND_605[5:0];
  _RAND_606 = {1{`RANDOM}};
  _T_3786_0 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  _T_3786_1 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  _T_3787_0 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  _T_3787_1 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  _T_3790 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  _T_3794 = _RAND_611[5:0];
  _RAND_612 = {1{`RANDOM}};
  _T_3795_0 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  _T_3795_1 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  _T_3796_0 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  _T_3796_1 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  _T_3799 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  _T_3803 = _RAND_617[5:0];
  _RAND_618 = {1{`RANDOM}};
  _T_3805_0 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  _T_3805_1 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  _T_3808 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  _T_3812 = _RAND_621[5:0];
  _RAND_622 = {1{`RANDOM}};
  _T_3814_0 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  _T_3814_1 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  _T_3817 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  _T_3821 = _RAND_625[5:0];
  _RAND_626 = {1{`RANDOM}};
  _T_3823_0 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  _T_3823_1 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  _T_3826 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  _T_3830 = _RAND_629[5:0];
  _RAND_630 = {1{`RANDOM}};
  _T_3832_0 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  _T_3832_1 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  _T_3835 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  _T_3839 = _RAND_633[5:0];
  _RAND_634 = {1{`RANDOM}};
  _T_3841_0 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  _T_3841_1 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  _T_3844 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  _T_3848 = _RAND_637[5:0];
  _RAND_638 = {1{`RANDOM}};
  _T_3850_0 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  _T_3850_1 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  _T_3853 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  _T_3857 = _RAND_641[5:0];
  _RAND_642 = {1{`RANDOM}};
  _T_3859_0 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  _T_3859_1 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  _T_3862 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  _T_3866 = _RAND_645[5:0];
  _RAND_646 = {1{`RANDOM}};
  _T_3867_0 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  _T_3867_1 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  _T_3868_0 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  _T_3868_1 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  _T_3871 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  _T_3875 = _RAND_651[5:0];
  _RAND_652 = {1{`RANDOM}};
  _T_3876_0 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  _T_3876_1 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  _T_3877_0 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  _T_3877_1 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  _T_3880 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  _T_3884 = _RAND_657[5:0];
  _RAND_658 = {1{`RANDOM}};
  _T_3885_0 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  _T_3885_1 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  _T_3886_0 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  _T_3886_1 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  _T_3889 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  _T_3893 = _RAND_663[5:0];
  _RAND_664 = {1{`RANDOM}};
  _T_3894_0 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  _T_3894_1 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  _T_3895_0 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  _T_3895_1 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  _T_3898 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  _T_3902 = _RAND_669[5:0];
  _RAND_670 = {1{`RANDOM}};
  _T_3903_0 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  _T_3903_1 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  _T_3904_0 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  _T_3904_1 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  _T_3907 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  _T_3911 = _RAND_675[5:0];
  _RAND_676 = {1{`RANDOM}};
  _T_3912_0 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  _T_3912_1 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  _T_3913_0 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  _T_3913_1 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  _T_3916 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  _T_3920 = _RAND_681[5:0];
  _RAND_682 = {1{`RANDOM}};
  _T_3921_0 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  _T_3921_1 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  _T_3922_0 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  _T_3922_1 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  _T_3925 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  _T_3929 = _RAND_687[5:0];
  _RAND_688 = {1{`RANDOM}};
  _T_3930_0 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  _T_3930_1 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  _T_3931_0 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  _T_3931_1 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  _T_3934 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  _T_3938 = _RAND_693[5:0];
  _RAND_694 = {1{`RANDOM}};
  _T_3939_0 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  _T_3939_1 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  _T_3940_0 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  _T_3940_1 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  _T_3943 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  _T_3947 = _RAND_699[5:0];
  _RAND_700 = {1{`RANDOM}};
  _T_3948_0 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  _T_3948_1 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  _T_3949_0 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  _T_3949_1 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  _T_3952 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  _T_3956 = _RAND_705[5:0];
  _RAND_706 = {1{`RANDOM}};
  _T_3957_0 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  _T_3957_1 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  _T_3958_0 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  _T_3958_1 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  _T_3961 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  _T_3965 = _RAND_711[5:0];
  _RAND_712 = {1{`RANDOM}};
  _T_3967_0 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  _T_3967_1 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  _T_3970 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  _T_3974 = _RAND_715[5:0];
  _RAND_716 = {1{`RANDOM}};
  _T_3976_0 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  _T_3976_1 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  _T_3979 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  _T_3983 = _RAND_719[5:0];
  _RAND_720 = {1{`RANDOM}};
  _T_3985_0 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  _T_3985_1 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  _T_3988 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  _T_3992 = _RAND_723[5:0];
  _RAND_724 = {1{`RANDOM}};
  _T_3993_0 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  _T_3993_1 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  _T_3994_0 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  _T_3994_1 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  _T_3997 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  _T_4001 = _RAND_729[5:0];
  _RAND_730 = {1{`RANDOM}};
  _T_4002_0 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  _T_4002_1 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  _T_4003_0 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  _T_4003_1 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  _T_4006 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  _T_4010 = _RAND_735[5:0];
  _RAND_736 = {1{`RANDOM}};
  _T_4011_0 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  _T_4011_1 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  _T_4012_0 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  _T_4012_1 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  _T_4015 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  _T_4019 = _RAND_741[5:0];
  _RAND_742 = {1{`RANDOM}};
  _T_4021_0 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  _T_4021_1 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  _T_4024 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  _T_4028 = _RAND_745[5:0];
  _RAND_746 = {1{`RANDOM}};
  _T_4030_0 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  _T_4030_1 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  _T_4033 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  _T_4037 = _RAND_749[5:0];
  _RAND_750 = {1{`RANDOM}};
  _T_4039_0 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  _T_4039_1 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  _T_4042 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  _T_4046 = _RAND_753[5:0];
  _RAND_754 = {1{`RANDOM}};
  _T_4047_0 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  _T_4047_1 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  _T_4048_0 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  _T_4048_1 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  _T_4051 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  _T_4055 = _RAND_759[5:0];
  _RAND_760 = {1{`RANDOM}};
  _T_4056_0 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  _T_4056_1 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  _T_4057_0 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  _T_4057_1 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  _T_4060 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  _T_4064 = _RAND_765[5:0];
  _RAND_766 = {1{`RANDOM}};
  _T_4065_0 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  _T_4065_1 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  _T_4066_0 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  _T_4066_1 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  _T_4069 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  _T_4073 = _RAND_771[5:0];
  _RAND_772 = {1{`RANDOM}};
  _T_4074_0 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  _T_4074_1 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  _T_4075_0 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  _T_4075_1 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  _T_4078 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  _T_4082 = _RAND_777[5:0];
  _RAND_778 = {1{`RANDOM}};
  _T_4083_0 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  _T_4083_1 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  _T_4084_0 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  _T_4084_1 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  _T_4087 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  _T_4091 = _RAND_783[5:0];
  _RAND_784 = {1{`RANDOM}};
  _T_4092_0 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  _T_4092_1 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  _T_4093_0 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  _T_4093_1 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  _T_4096 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  _T_4100 = _RAND_789[5:0];
  _RAND_790 = {1{`RANDOM}};
  _T_4102_0 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  _T_4102_1 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  _T_4105 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  _T_4109 = _RAND_793[5:0];
  _RAND_794 = {1{`RANDOM}};
  _T_4111_0 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  _T_4111_1 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  _T_4114 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  _T_4118 = _RAND_797[5:0];
  _RAND_798 = {1{`RANDOM}};
  _T_4120_0 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  _T_4120_1 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  _T_4123 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  _T_4127 = _RAND_801[5:0];
  _RAND_802 = {1{`RANDOM}};
  _T_4128_0 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  _T_4128_1 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  _T_4129_0 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  _T_4129_1 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  _T_4132 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  _T_4136 = _RAND_807[5:0];
  _RAND_808 = {1{`RANDOM}};
  _T_4137_0 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  _T_4137_1 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  _T_4138_0 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  _T_4138_1 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  _T_4141 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  _T_4145 = _RAND_813[5:0];
  _RAND_814 = {1{`RANDOM}};
  _T_4146_0 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  _T_4146_1 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  _T_4147_0 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  _T_4147_1 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  _T_4150 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  _T_4154 = _RAND_819[5:0];
  _RAND_820 = {1{`RANDOM}};
  _T_4156_0 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  _T_4156_1 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  _T_4159 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  _T_4163 = _RAND_823[5:0];
  _RAND_824 = {1{`RANDOM}};
  _T_4165_0 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  _T_4165_1 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  _T_4168 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  _T_4172 = _RAND_827[5:0];
  _RAND_828 = {1{`RANDOM}};
  _T_4174_0 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  _T_4174_1 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  _T_4177 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  _T_4181 = _RAND_831[5:0];
  _RAND_832 = {1{`RANDOM}};
  _T_4183_0 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  _T_4183_1 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  _T_4186 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  _T_4190 = _RAND_835[5:0];
  _RAND_836 = {1{`RANDOM}};
  _T_4192_0 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  _T_4192_1 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  _T_4195 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  _T_4199 = _RAND_839[5:0];
  _RAND_840 = {1{`RANDOM}};
  _T_4201_0 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  _T_4201_1 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  _T_4204 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  _T_4208 = _RAND_843[5:0];
  _RAND_844 = {1{`RANDOM}};
  _T_4210_0 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  _T_4210_1 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  _T_4213 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  _T_4217 = _RAND_847[5:0];
  _RAND_848 = {1{`RANDOM}};
  _T_4219_0 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  _T_4219_1 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  _T_4222 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  _T_4226 = _RAND_851[5:0];
  _RAND_852 = {1{`RANDOM}};
  _T_4228_0 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  _T_4228_1 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  _T_4231 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  _T_4235 = _RAND_855[5:0];
  _RAND_856 = {1{`RANDOM}};
  _T_4237_0 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  _T_4237_1 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  _T_4240 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  _T_4244 = _RAND_859[5:0];
  _RAND_860 = {1{`RANDOM}};
  _T_4246_0 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  _T_4246_1 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  _T_4249 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  _T_4253 = _RAND_863[5:0];
  _RAND_864 = {1{`RANDOM}};
  _T_4255_0 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  _T_4255_1 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  _T_4258 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  _T_4262 = _RAND_867[5:0];
  _RAND_868 = {1{`RANDOM}};
  _T_4264_0 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  _T_4264_1 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  _T_4267 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  _T_4271 = _RAND_871[5:0];
  _RAND_872 = {1{`RANDOM}};
  _T_4273_0 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  _T_4273_1 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  _T_4276 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  _T_4280 = _RAND_875[5:0];
  _RAND_876 = {1{`RANDOM}};
  _T_4282_0 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  _T_4282_1 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  _T_4285 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  _T_4289 = _RAND_879[5:0];
  _RAND_880 = {1{`RANDOM}};
  _T_4291_0 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  _T_4291_1 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  _T_4294 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  _T_4298 = _RAND_883[5:0];
  _RAND_884 = {1{`RANDOM}};
  _T_4300_0 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  _T_4300_1 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  _T_4303 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  _T_4307 = _RAND_887[5:0];
  _RAND_888 = {1{`RANDOM}};
  _T_4309_0 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  _T_4309_1 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  _T_4312 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  _T_4316 = _RAND_891[5:0];
  _RAND_892 = {1{`RANDOM}};
  _T_4318_0 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  _T_4318_1 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  _T_4321 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  _T_4325 = _RAND_895[5:0];
  _RAND_896 = {1{`RANDOM}};
  _T_4327_0 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  _T_4327_1 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  _T_4330 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  _T_4334 = _RAND_899[5:0];
  _RAND_900 = {1{`RANDOM}};
  _T_4336_0 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  _T_4336_1 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  _T_4339 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  _T_4343 = _RAND_903[5:0];
  _RAND_904 = {1{`RANDOM}};
  _T_4345_0 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  _T_4345_1 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  _T_4348 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  _T_4352 = _RAND_907[5:0];
  _RAND_908 = {1{`RANDOM}};
  _T_4354_0 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  _T_4354_1 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  _T_4357 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  _T_4361 = _RAND_911[5:0];
  _RAND_912 = {1{`RANDOM}};
  _T_4363_0 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  _T_4363_1 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  _T_4366 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  _T_4370 = _RAND_915[5:0];
  _RAND_916 = {1{`RANDOM}};
  _T_4372_0 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  _T_4372_1 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  _T_4375 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  _T_4379 = _RAND_919[5:0];
  _RAND_920 = {1{`RANDOM}};
  _T_4381_0 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  _T_4381_1 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  _T_4384 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  _T_4388 = _RAND_923[5:0];
  _RAND_924 = {1{`RANDOM}};
  _T_4390_0 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  _T_4390_1 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  _T_4393 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  _T_4397 = _RAND_927[5:0];
  _RAND_928 = {1{`RANDOM}};
  _T_4399_0 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  _T_4399_1 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  _T_4402 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  _T_4406 = _RAND_931[5:0];
  _RAND_932 = {1{`RANDOM}};
  _T_4408_0 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  _T_4408_1 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  _T_4411 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  _T_4415 = _RAND_935[5:0];
  _RAND_936 = {1{`RANDOM}};
  _T_4417_0 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  _T_4417_1 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  _T_4420 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  _T_4424 = _RAND_939[5:0];
  _RAND_940 = {1{`RANDOM}};
  _T_4426_0 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  _T_4426_1 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  _T_4429 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  _T_4433 = _RAND_943[5:0];
  _RAND_944 = {1{`RANDOM}};
  _T_4435_0 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  _T_4435_1 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  _T_4438 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  _T_4442 = _RAND_947[5:0];
  _RAND_948 = {1{`RANDOM}};
  _T_4444_0 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  _T_4444_1 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  _T_4447 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  _T_4451 = _RAND_951[5:0];
  _RAND_952 = {1{`RANDOM}};
  _T_4453_0 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  _T_4453_1 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  _T_4456 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  _T_4460 = _RAND_955[5:0];
  _RAND_956 = {1{`RANDOM}};
  _T_4462_0 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  _T_4462_1 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  _T_4465 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  _T_4469 = _RAND_959[5:0];
  _RAND_960 = {1{`RANDOM}};
  _T_4471_0 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  _T_4471_1 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  _T_4474 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  _T_4478 = _RAND_963[5:0];
  _RAND_964 = {1{`RANDOM}};
  _T_4480_0 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  _T_4480_1 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  _T_4483 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  _T_4487 = _RAND_967[5:0];
  _RAND_968 = {1{`RANDOM}};
  _T_4489_0 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  _T_4489_1 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  _T_4492 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  _T_4496 = _RAND_971[5:0];
  _RAND_972 = {1{`RANDOM}};
  _T_4498_0 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  _T_4498_1 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  _T_4501 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  _T_4505 = _RAND_975[5:0];
  _RAND_976 = {1{`RANDOM}};
  _T_4507_0 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  _T_4507_1 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  _T_4510 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  _T_4514 = _RAND_979[5:0];
  _RAND_980 = {1{`RANDOM}};
  _T_4516_0 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  _T_4516_1 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  _T_4519 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  _T_4523 = _RAND_983[5:0];
  _RAND_984 = {1{`RANDOM}};
  _T_4525_0 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  _T_4525_1 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  _T_4528 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  _T_4532 = _RAND_987[5:0];
  _RAND_988 = {1{`RANDOM}};
  _T_4534_0 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  _T_4534_1 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  _T_4537 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  _T_4541 = _RAND_991[5:0];
  _RAND_992 = {1{`RANDOM}};
  _T_4543_0 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  _T_4543_1 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  _T_4546 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  _T_4550 = _RAND_995[5:0];
  _RAND_996 = {1{`RANDOM}};
  _T_4552_0 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  _T_4552_1 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  _T_4555 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  _T_4559 = _RAND_999[5:0];
  _RAND_1000 = {1{`RANDOM}};
  _T_4561_0 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  _T_4561_1 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  _T_4564 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  _T_4568 = _RAND_1003[5:0];
  _RAND_1004 = {1{`RANDOM}};
  _T_4570_0 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  _T_4570_1 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  _T_4573 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  _T_4577 = _RAND_1007[5:0];
  _RAND_1008 = {1{`RANDOM}};
  _T_4579_0 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  _T_4579_1 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  _T_4582 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  _T_4586 = _RAND_1011[5:0];
  _RAND_1012 = {1{`RANDOM}};
  _T_4588_0 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  _T_4588_1 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  _T_4591 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  _T_4595 = _RAND_1015[5:0];
  _RAND_1016 = {1{`RANDOM}};
  _T_4597_0 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  _T_4597_1 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  _T_4600 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  _T_4604 = _RAND_1019[5:0];
  _RAND_1020 = {1{`RANDOM}};
  _T_4606_0 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  _T_4606_1 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  _T_4609 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  _T_4613 = _RAND_1023[5:0];
  _RAND_1024 = {1{`RANDOM}};
  _T_4615_0 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  _T_4615_1 = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  _T_4618 = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  _T_4622 = _RAND_1027[5:0];
  _RAND_1028 = {1{`RANDOM}};
  _T_4624_0 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  _T_4624_1 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  _T_4627 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  _T_4631 = _RAND_1031[5:0];
  _RAND_1032 = {1{`RANDOM}};
  _T_4633_0 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  _T_4633_1 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  _T_4636 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  _T_4640 = _RAND_1035[5:0];
  _RAND_1036 = {1{`RANDOM}};
  _T_4642_0 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  _T_4642_1 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  _T_4645 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  pixelColorSprite = _RAND_1039[5:0];
  _RAND_1040 = {1{`RANDOM}};
  pixelColorSpriteValid = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  _T_4648_0 = _RAND_1041[0:0];
  _RAND_1042 = {1{`RANDOM}};
  _T_4648_1 = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  _T_4648_2 = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  _T_4655 = _RAND_1044[3:0];
  _RAND_1045 = {1{`RANDOM}};
  _T_4656 = _RAND_1045[3:0];
  _RAND_1046 = {1{`RANDOM}};
  _T_4657 = _RAND_1046[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ScaleCounterReg <= 2'h0;
    end else if (run) begin
      if (_T) begin
        ScaleCounterReg <= 2'h0;
      end else begin
        ScaleCounterReg <= _T_8;
      end
    end
    if (reset) begin
      CounterXReg <= 10'h0;
    end else if (run) begin
      if (_T) begin
        if (_T_1) begin
          CounterXReg <= 10'h0;
        end else begin
          CounterXReg <= _T_6;
        end
      end
    end
    if (reset) begin
      CounterYReg <= 10'h0;
    end else if (run) begin
      if (_T) begin
        if (_T_1) begin
          if (_T_2) begin
            CounterYReg <= 10'h0;
          end else begin
            CounterYReg <= _T_4;
          end
        end
      end
    end
    if (reset) begin
      backMemoryRestoreCounter <= 12'h0;
    end else if (restoreEnabled) begin
      backMemoryRestoreCounter <= _T_370;
    end
    _T_14_0 <= _T_14_1;
    _T_14_1 <= _T_14_2;
    _T_14_2 <= _T_14_3;
    _T_14_3 <= ~Hsync;
    _T_16_0 <= _T_16_1;
    _T_16_1 <= _T_16_2;
    _T_16_2 <= _T_16_3;
    _T_16_3 <= ~Vsync;
    if (reset) begin
      frameClockCount <= 21'h0;
    end else if (_T_19) begin
      frameClockCount <= 21'h0;
    end else begin
      frameClockCount <= _T_21;
    end
    if (reset) begin
      spriteXPositionReg_0 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_0 <= io_spriteXPosition_0;
    end
    if (reset) begin
      spriteXPositionReg_1 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_1 <= io_spriteXPosition_1;
    end
    if (reset) begin
      spriteXPositionReg_2 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_2 <= io_spriteXPosition_2;
    end
    if (reset) begin
      spriteXPositionReg_3 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_3 <= io_spriteXPosition_3;
    end
    if (reset) begin
      spriteXPositionReg_4 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_4 <= io_spriteXPosition_4;
    end
    if (reset) begin
      spriteXPositionReg_5 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_5 <= io_spriteXPosition_5;
    end
    if (reset) begin
      spriteXPositionReg_6 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_6 <= io_spriteXPosition_6;
    end
    if (reset) begin
      spriteXPositionReg_7 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_7 <= io_spriteXPosition_7;
    end
    if (reset) begin
      spriteXPositionReg_8 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_8 <= io_spriteXPosition_8;
    end
    if (reset) begin
      spriteXPositionReg_9 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_9 <= io_spriteXPosition_9;
    end
    if (reset) begin
      spriteXPositionReg_10 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_10 <= io_spriteXPosition_10;
    end
    if (reset) begin
      spriteXPositionReg_11 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_11 <= io_spriteXPosition_11;
    end
    if (reset) begin
      spriteXPositionReg_12 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_12 <= io_spriteXPosition_12;
    end
    if (reset) begin
      spriteXPositionReg_13 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_13 <= io_spriteXPosition_13;
    end
    if (reset) begin
      spriteXPositionReg_14 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_14 <= io_spriteXPosition_14;
    end
    if (reset) begin
      spriteXPositionReg_15 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_15 <= io_spriteXPosition_15;
    end
    if (reset) begin
      spriteXPositionReg_16 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_16 <= io_spriteXPosition_16;
    end
    if (reset) begin
      spriteXPositionReg_17 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_17 <= io_spriteXPosition_17;
    end
    if (reset) begin
      spriteXPositionReg_18 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_18 <= io_spriteXPosition_18;
    end
    if (reset) begin
      spriteXPositionReg_19 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_19 <= io_spriteXPosition_19;
    end
    if (reset) begin
      spriteXPositionReg_20 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_20 <= io_spriteXPosition_20;
    end
    if (reset) begin
      spriteXPositionReg_21 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_21 <= io_spriteXPosition_21;
    end
    if (reset) begin
      spriteXPositionReg_22 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_22 <= io_spriteXPosition_22;
    end
    if (reset) begin
      spriteXPositionReg_23 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_23 <= io_spriteXPosition_23;
    end
    if (reset) begin
      spriteXPositionReg_24 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_24 <= io_spriteXPosition_24;
    end
    if (reset) begin
      spriteXPositionReg_25 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_25 <= io_spriteXPosition_25;
    end
    if (reset) begin
      spriteXPositionReg_26 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_26 <= io_spriteXPosition_26;
    end
    if (reset) begin
      spriteXPositionReg_27 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_27 <= io_spriteXPosition_27;
    end
    if (reset) begin
      spriteXPositionReg_28 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_28 <= io_spriteXPosition_28;
    end
    if (reset) begin
      spriteXPositionReg_29 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_29 <= io_spriteXPosition_29;
    end
    if (reset) begin
      spriteXPositionReg_30 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_30 <= io_spriteXPosition_30;
    end
    if (reset) begin
      spriteXPositionReg_31 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_31 <= io_spriteXPosition_31;
    end
    if (reset) begin
      spriteXPositionReg_32 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_32 <= io_spriteXPosition_32;
    end
    if (reset) begin
      spriteXPositionReg_33 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_33 <= io_spriteXPosition_33;
    end
    if (reset) begin
      spriteXPositionReg_34 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_34 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_35 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_35 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_36 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_36 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_37 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_37 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_38 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_38 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_39 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_39 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_40 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_40 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_41 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_41 <= io_spriteXPosition_41;
    end
    if (reset) begin
      spriteXPositionReg_42 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_42 <= io_spriteXPosition_42;
    end
    if (reset) begin
      spriteXPositionReg_43 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_43 <= io_spriteXPosition_43;
    end
    if (reset) begin
      spriteXPositionReg_44 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_44 <= io_spriteXPosition_44;
    end
    if (reset) begin
      spriteXPositionReg_45 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_45 <= io_spriteXPosition_45;
    end
    if (reset) begin
      spriteXPositionReg_46 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_46 <= io_spriteXPosition_46;
    end
    if (reset) begin
      spriteXPositionReg_47 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_47 <= io_spriteXPosition_47;
    end
    if (reset) begin
      spriteXPositionReg_48 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_48 <= io_spriteXPosition_48;
    end
    if (reset) begin
      spriteXPositionReg_49 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_49 <= io_spriteXPosition_49;
    end
    if (reset) begin
      spriteXPositionReg_50 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_50 <= io_spriteXPosition_50;
    end
    if (reset) begin
      spriteXPositionReg_51 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_51 <= io_spriteXPosition_51;
    end
    if (reset) begin
      spriteXPositionReg_52 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_52 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_53 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_53 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_54 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_54 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_55 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_55 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_56 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_56 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_57 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_57 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_58 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_58 <= 11'sh1e0;
    end
    if (reset) begin
      spriteXPositionReg_59 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_59 <= 11'sh200;
    end
    if (reset) begin
      spriteXPositionReg_60 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_60 <= 11'sh220;
    end
    if (reset) begin
      spriteXPositionReg_61 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_61 <= 11'sh1e0;
    end
    if (reset) begin
      spriteXPositionReg_62 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_62 <= 11'sh200;
    end
    if (reset) begin
      spriteXPositionReg_63 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_63 <= 11'sh220;
    end
    if (reset) begin
      spriteXPositionReg_64 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_64 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_65 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_65 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_66 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_66 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_67 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_67 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_68 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_68 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_69 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_69 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_70 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_70 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_71 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_71 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_72 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_72 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_73 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_73 <= 11'sh140;
    end
    if (reset) begin
      spriteXPositionReg_74 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_74 <= 11'sh120;
    end
    if (reset) begin
      spriteXPositionReg_75 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_75 <= 11'sh100;
    end
    if (reset) begin
      spriteXPositionReg_76 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_76 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_77 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_77 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_78 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_78 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_79 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_79 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_80 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_80 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_81 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_81 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_82 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_82 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_83 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_83 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_84 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_84 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_85 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_85 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_86 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_86 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_87 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_87 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_88 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_88 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_89 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_89 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_90 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_90 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_91 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_91 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_92 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_92 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_93 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_93 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_94 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_94 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_95 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_95 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_96 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_96 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_97 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_97 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_98 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_98 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_99 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_99 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_100 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_100 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_101 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_101 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_102 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_102 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_103 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_103 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_104 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_104 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_105 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_105 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_106 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_106 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_107 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_107 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_108 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_108 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_109 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_109 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_110 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_110 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_111 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_111 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_112 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_112 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_113 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_113 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_114 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_114 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_115 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_115 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_116 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_116 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_117 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_117 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_118 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_118 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_119 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_119 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_120 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_120 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_121 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_121 <= 11'sh2bc;
    end
    if (reset) begin
      spriteXPositionReg_122 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_122 <= io_spriteXPosition_122;
    end
    if (reset) begin
      spriteXPositionReg_123 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_123 <= io_spriteXPosition_123;
    end
    if (reset) begin
      spriteXPositionReg_124 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_124 <= io_spriteXPosition_124;
    end
    if (reset) begin
      spriteXPositionReg_125 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_125 <= io_spriteXPosition_125;
    end
    if (reset) begin
      spriteXPositionReg_126 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_126 <= io_spriteXPosition_126;
    end
    if (reset) begin
      spriteXPositionReg_127 <= 11'sh0;
    end else if (io_newFrame) begin
      spriteXPositionReg_127 <= io_spriteXPosition_127;
    end
    if (reset) begin
      spriteYPositionReg_0 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_0 <= io_spriteYPosition_0;
    end
    if (reset) begin
      spriteYPositionReg_1 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_1 <= io_spriteYPosition_1;
    end
    if (reset) begin
      spriteYPositionReg_2 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_2 <= io_spriteYPosition_2;
    end
    if (reset) begin
      spriteYPositionReg_3 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_3 <= io_spriteYPosition_3;
    end
    if (reset) begin
      spriteYPositionReg_4 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_4 <= io_spriteYPosition_4;
    end
    if (reset) begin
      spriteYPositionReg_5 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_5 <= io_spriteYPosition_5;
    end
    if (reset) begin
      spriteYPositionReg_6 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_6 <= io_spriteYPosition_6;
    end
    if (reset) begin
      spriteYPositionReg_7 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_7 <= io_spriteYPosition_7;
    end
    if (reset) begin
      spriteYPositionReg_8 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_8 <= io_spriteYPosition_8;
    end
    if (reset) begin
      spriteYPositionReg_9 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_9 <= io_spriteYPosition_9;
    end
    if (reset) begin
      spriteYPositionReg_10 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_10 <= io_spriteYPosition_10;
    end
    if (reset) begin
      spriteYPositionReg_11 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_11 <= io_spriteYPosition_11;
    end
    if (reset) begin
      spriteYPositionReg_12 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_12 <= io_spriteYPosition_12;
    end
    if (reset) begin
      spriteYPositionReg_13 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_13 <= io_spriteYPosition_13;
    end
    if (reset) begin
      spriteYPositionReg_14 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_14 <= io_spriteYPosition_14;
    end
    if (reset) begin
      spriteYPositionReg_15 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_15 <= io_spriteYPosition_15;
    end
    if (reset) begin
      spriteYPositionReg_16 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_16 <= io_spriteYPosition_16;
    end
    if (reset) begin
      spriteYPositionReg_17 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_17 <= io_spriteYPosition_17;
    end
    if (reset) begin
      spriteYPositionReg_18 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_18 <= io_spriteYPosition_18;
    end
    if (reset) begin
      spriteYPositionReg_19 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_19 <= io_spriteYPosition_19;
    end
    if (reset) begin
      spriteYPositionReg_20 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_20 <= io_spriteYPosition_20;
    end
    if (reset) begin
      spriteYPositionReg_21 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_21 <= io_spriteYPosition_21;
    end
    if (reset) begin
      spriteYPositionReg_22 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_22 <= io_spriteYPosition_22;
    end
    if (reset) begin
      spriteYPositionReg_23 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_23 <= io_spriteYPosition_23;
    end
    if (reset) begin
      spriteYPositionReg_24 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_24 <= io_spriteYPosition_24;
    end
    if (reset) begin
      spriteYPositionReg_25 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_25 <= io_spriteYPosition_25;
    end
    if (reset) begin
      spriteYPositionReg_26 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_26 <= io_spriteYPosition_26;
    end
    if (reset) begin
      spriteYPositionReg_27 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_27 <= io_spriteYPosition_27;
    end
    if (reset) begin
      spriteYPositionReg_28 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_28 <= io_spriteYPosition_28;
    end
    if (reset) begin
      spriteYPositionReg_29 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_29 <= io_spriteYPosition_29;
    end
    if (reset) begin
      spriteYPositionReg_30 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_30 <= io_spriteYPosition_30;
    end
    if (reset) begin
      spriteYPositionReg_31 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_31 <= io_spriteYPosition_31;
    end
    if (reset) begin
      spriteYPositionReg_32 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_32 <= io_spriteYPosition_32;
    end
    if (reset) begin
      spriteYPositionReg_33 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_33 <= io_spriteYPosition_33;
    end
    if (reset) begin
      spriteYPositionReg_34 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_34 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_35 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_35 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_36 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_36 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_37 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_37 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_38 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_38 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_39 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_39 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_40 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_40 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_41 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_41 <= io_spriteYPosition_41;
    end
    if (reset) begin
      spriteYPositionReg_42 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_42 <= io_spriteYPosition_42;
    end
    if (reset) begin
      spriteYPositionReg_43 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_43 <= io_spriteYPosition_43;
    end
    if (reset) begin
      spriteYPositionReg_44 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_44 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_45 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_45 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_46 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_46 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_47 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_47 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_48 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_48 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_49 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_49 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_50 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_50 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_51 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_51 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_52 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_52 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_53 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_53 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_54 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_54 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_55 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_55 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_56 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_56 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_57 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_57 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_58 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_58 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_59 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_59 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_60 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_60 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_61 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_61 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_62 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_62 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_63 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_63 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_70 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_70 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_71 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_71 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_72 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_72 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_73 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_73 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_74 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_74 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_75 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_75 <= 10'sh40;
    end
    if (reset) begin
      spriteYPositionReg_76 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_76 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_77 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_77 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_78 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_78 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_79 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_79 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_80 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_80 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_81 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_81 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_82 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_82 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_83 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_83 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_84 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_84 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_85 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_85 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_86 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_86 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_87 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_87 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_88 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_88 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_89 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_89 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_90 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_90 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_91 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_91 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_92 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_92 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_93 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_93 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_94 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_94 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_95 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_95 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_96 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_96 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_97 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_97 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_98 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_98 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_99 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_99 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_100 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_100 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_101 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_101 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_102 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_102 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_103 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_103 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_104 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_104 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_105 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_105 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_106 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_106 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_107 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_107 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_108 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_108 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_109 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_109 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_110 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_110 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_111 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_111 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_112 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_112 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_113 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_113 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_114 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_114 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_115 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_115 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_116 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_116 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_117 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_117 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_118 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_118 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_119 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_119 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_120 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_120 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_121 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_121 <= 10'sh20;
    end
    if (reset) begin
      spriteYPositionReg_122 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_122 <= io_spriteYPosition_122;
    end
    if (reset) begin
      spriteYPositionReg_123 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_123 <= io_spriteYPosition_123;
    end
    if (reset) begin
      spriteYPositionReg_124 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_124 <= io_spriteYPosition_124;
    end
    if (reset) begin
      spriteYPositionReg_125 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_125 <= io_spriteYPosition_125;
    end
    if (reset) begin
      spriteYPositionReg_126 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_126 <= io_spriteYPosition_126;
    end
    if (reset) begin
      spriteYPositionReg_127 <= 10'sh0;
    end else if (io_newFrame) begin
      spriteYPositionReg_127 <= io_spriteYPosition_127;
    end
    spriteVisibleReg_0 <= reset | _GEN_269;
    spriteVisibleReg_1 <= reset | _GEN_270;
    spriteVisibleReg_2 <= reset | _GEN_271;
    spriteVisibleReg_3 <= reset | _GEN_272;
    spriteVisibleReg_4 <= reset | _GEN_273;
    spriteVisibleReg_5 <= reset | _GEN_274;
    spriteVisibleReg_6 <= reset | _GEN_275;
    spriteVisibleReg_7 <= reset | _GEN_276;
    spriteVisibleReg_8 <= reset | _GEN_277;
    spriteVisibleReg_9 <= reset | _GEN_278;
    spriteVisibleReg_10 <= reset | _GEN_279;
    spriteVisibleReg_11 <= reset | _GEN_280;
    spriteVisibleReg_12 <= reset | _GEN_281;
    spriteVisibleReg_13 <= reset | _GEN_282;
    spriteVisibleReg_14 <= reset | _GEN_283;
    spriteVisibleReg_15 <= reset | _GEN_284;
    spriteVisibleReg_16 <= reset | _GEN_285;
    spriteVisibleReg_17 <= reset | _GEN_286;
    spriteVisibleReg_18 <= reset | _GEN_287;
    spriteVisibleReg_19 <= reset | _GEN_288;
    spriteVisibleReg_20 <= reset | _GEN_289;
    spriteVisibleReg_21 <= reset | _GEN_290;
    spriteVisibleReg_22 <= reset | _GEN_291;
    spriteVisibleReg_23 <= reset | _GEN_292;
    spriteVisibleReg_24 <= reset | _GEN_293;
    spriteVisibleReg_25 <= reset | _GEN_294;
    spriteVisibleReg_26 <= reset | _GEN_295;
    spriteVisibleReg_27 <= reset | _GEN_296;
    spriteVisibleReg_28 <= reset | _GEN_297;
    spriteVisibleReg_29 <= reset | _GEN_298;
    spriteVisibleReg_30 <= reset | _GEN_299;
    spriteVisibleReg_31 <= reset | _GEN_300;
    spriteVisibleReg_32 <= reset | _GEN_301;
    spriteVisibleReg_33 <= reset | _GEN_302;
    spriteVisibleReg_41 <= reset | _GEN_310;
    spriteVisibleReg_42 <= reset | _GEN_311;
    spriteVisibleReg_43 <= reset | _GEN_312;
    spriteVisibleReg_44 <= reset | _GEN_313;
    spriteVisibleReg_45 <= reset | _GEN_314;
    spriteVisibleReg_46 <= reset | _GEN_315;
    spriteVisibleReg_47 <= reset | _GEN_316;
    spriteVisibleReg_48 <= reset | _GEN_317;
    spriteVisibleReg_49 <= reset | _GEN_318;
    spriteVisibleReg_50 <= reset | _GEN_319;
    spriteVisibleReg_51 <= reset | _GEN_320;
    spriteVisibleReg_55 <= reset | _GEN_324;
    spriteVisibleReg_56 <= reset | _GEN_325;
    spriteVisibleReg_57 <= reset | _GEN_326;
    spriteVisibleReg_61 <= reset | _GEN_330;
    spriteVisibleReg_62 <= reset | _GEN_331;
    spriteVisibleReg_63 <= reset | _GEN_332;
    spriteVisibleReg_64 <= reset | _GEN_333;
    spriteVisibleReg_65 <= reset | _GEN_334;
    spriteVisibleReg_66 <= reset | _GEN_335;
    spriteVisibleReg_70 <= reset | _GEN_339;
    spriteVisibleReg_71 <= reset | _GEN_340;
    spriteVisibleReg_72 <= reset | _GEN_341;
    if (reset) begin
      spriteFlipVerticalReg_122 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_122 <= io_spriteFlipVertical_122;
    end
    if (reset) begin
      spriteFlipVerticalReg_123 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_123 <= io_spriteFlipVertical_123;
    end
    if (reset) begin
      spriteFlipVerticalReg_124 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_124 <= io_spriteFlipVertical_124;
    end
    if (reset) begin
      spriteFlipVerticalReg_125 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_125 <= io_spriteFlipVertical_125;
    end
    if (reset) begin
      spriteFlipVerticalReg_126 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_126 <= io_spriteFlipVertical_126;
    end
    if (reset) begin
      spriteFlipVerticalReg_127 <= 1'h0;
    end else if (io_newFrame) begin
      spriteFlipVerticalReg_127 <= io_spriteFlipVertical_127;
    end
    if (reset) begin
      viewBoxXReg_0 <= 10'h0;
    end else if (io_newFrame) begin
      viewBoxXReg_0 <= io_viewBoxX_0;
    end
    if (reset) begin
      missingFrameErrorReg <= 1'h0;
    end else begin
      missingFrameErrorReg <= _GEN_660;
    end
    if (reset) begin
      backBufferWriteErrorReg <= 1'h0;
    end else if (_T_411) begin
      backBufferWriteErrorReg <= _GEN_668;
    end
    if (reset) begin
      viewBoxOutOfRangeErrorReg <= 1'h0;
    end else begin
      viewBoxOutOfRangeErrorReg <= _GEN_657;
    end
    if (reset) begin
      newFrameStikyReg <= 1'h0;
    end else if (_T_43) begin
      newFrameStikyReg <= 1'h0;
    end else begin
      newFrameStikyReg <= _GEN_658;
    end
    _T_43 <= io_frameUpdateDone;
    backTileMemoryDataRead_0_0 <= backTileMemories_0_0_io_dataRead;
    backTileMemoryDataRead_0_1 <= backTileMemories_0_1_io_dataRead;
    backTileMemoryDataRead_0_2 <= backTileMemories_0_2_io_dataRead;
    backTileMemoryDataRead_0_3 <= backTileMemories_0_3_io_dataRead;
    backTileMemoryDataRead_0_4 <= backTileMemories_0_4_io_dataRead;
    backTileMemoryDataRead_0_5 <= backTileMemories_0_5_io_dataRead;
    backTileMemoryDataRead_0_6 <= backTileMemories_0_6_io_dataRead;
    backTileMemoryDataRead_0_7 <= backTileMemories_0_7_io_dataRead;
    backTileMemoryDataRead_0_8 <= backTileMemories_0_8_io_dataRead;
    backTileMemoryDataRead_0_9 <= backTileMemories_0_9_io_dataRead;
    backTileMemoryDataRead_0_10 <= backTileMemories_0_10_io_dataRead;
    backTileMemoryDataRead_0_11 <= backTileMemories_0_11_io_dataRead;
    backTileMemoryDataRead_0_12 <= backTileMemories_0_12_io_dataRead;
    backTileMemoryDataRead_0_13 <= backTileMemories_0_13_io_dataRead;
    backTileMemoryDataRead_0_14 <= backTileMemories_0_14_io_dataRead;
    backTileMemoryDataRead_0_15 <= backTileMemories_0_15_io_dataRead;
    backTileMemoryDataRead_0_16 <= backTileMemories_0_16_io_dataRead;
    backTileMemoryDataRead_0_17 <= backTileMemories_0_17_io_dataRead;
    backTileMemoryDataRead_0_18 <= backTileMemories_0_18_io_dataRead;
    backTileMemoryDataRead_0_19 <= backTileMemories_0_19_io_dataRead;
    backTileMemoryDataRead_0_20 <= backTileMemories_0_20_io_dataRead;
    backTileMemoryDataRead_0_21 <= backTileMemories_0_21_io_dataRead;
    backTileMemoryDataRead_0_22 <= backTileMemories_0_22_io_dataRead;
    backTileMemoryDataRead_0_23 <= backTileMemories_0_23_io_dataRead;
    backTileMemoryDataRead_0_24 <= backTileMemories_0_24_io_dataRead;
    backTileMemoryDataRead_0_25 <= backTileMemories_0_25_io_dataRead;
    backTileMemoryDataRead_0_26 <= backTileMemories_0_26_io_dataRead;
    backTileMemoryDataRead_0_27 <= backTileMemories_0_27_io_dataRead;
    backTileMemoryDataRead_0_28 <= backTileMemories_0_28_io_dataRead;
    backTileMemoryDataRead_0_29 <= backTileMemories_0_29_io_dataRead;
    backTileMemoryDataRead_0_30 <= backTileMemories_0_30_io_dataRead;
    backTileMemoryDataRead_0_31 <= backTileMemories_0_31_io_dataRead;
    backTileMemoryDataRead_1_0 <= backTileMemories_1_0_io_dataRead;
    backTileMemoryDataRead_1_1 <= backTileMemories_1_1_io_dataRead;
    backTileMemoryDataRead_1_2 <= backTileMemories_1_2_io_dataRead;
    backTileMemoryDataRead_1_3 <= backTileMemories_1_3_io_dataRead;
    backTileMemoryDataRead_1_4 <= backTileMemories_1_4_io_dataRead;
    backTileMemoryDataRead_1_5 <= backTileMemories_1_5_io_dataRead;
    backTileMemoryDataRead_1_6 <= backTileMemories_1_6_io_dataRead;
    backTileMemoryDataRead_1_7 <= backTileMemories_1_7_io_dataRead;
    backTileMemoryDataRead_1_8 <= backTileMemories_1_8_io_dataRead;
    backTileMemoryDataRead_1_9 <= backTileMemories_1_9_io_dataRead;
    backTileMemoryDataRead_1_10 <= backTileMemories_1_10_io_dataRead;
    backTileMemoryDataRead_1_11 <= backTileMemories_1_11_io_dataRead;
    backTileMemoryDataRead_1_12 <= backTileMemories_1_12_io_dataRead;
    backTileMemoryDataRead_1_13 <= backTileMemories_1_13_io_dataRead;
    backTileMemoryDataRead_1_14 <= backTileMemories_1_14_io_dataRead;
    backTileMemoryDataRead_1_15 <= backTileMemories_1_15_io_dataRead;
    backTileMemoryDataRead_1_16 <= backTileMemories_1_16_io_dataRead;
    backTileMemoryDataRead_1_17 <= backTileMemories_1_17_io_dataRead;
    backTileMemoryDataRead_1_18 <= backTileMemories_1_18_io_dataRead;
    backTileMemoryDataRead_1_19 <= backTileMemories_1_19_io_dataRead;
    backTileMemoryDataRead_1_20 <= backTileMemories_1_20_io_dataRead;
    backTileMemoryDataRead_1_21 <= backTileMemories_1_21_io_dataRead;
    backTileMemoryDataRead_1_22 <= backTileMemories_1_22_io_dataRead;
    backTileMemoryDataRead_1_23 <= backTileMemories_1_23_io_dataRead;
    backTileMemoryDataRead_1_24 <= backTileMemories_1_24_io_dataRead;
    backTileMemoryDataRead_1_25 <= backTileMemories_1_25_io_dataRead;
    backTileMemoryDataRead_1_26 <= backTileMemories_1_26_io_dataRead;
    backTileMemoryDataRead_1_27 <= backTileMemories_1_27_io_dataRead;
    backTileMemoryDataRead_1_28 <= backTileMemories_1_28_io_dataRead;
    backTileMemoryDataRead_1_29 <= backTileMemories_1_29_io_dataRead;
    backTileMemoryDataRead_1_30 <= backTileMemories_1_30_io_dataRead;
    backTileMemoryDataRead_1_31 <= backTileMemories_1_31_io_dataRead;
    if (reset) begin
      backMemoryCopyCounter <= 12'h0;
    end else if (preDisplayArea) begin
      if (_T_365) begin
        backMemoryCopyCounter <= _T_367;
      end
    end else begin
      backMemoryCopyCounter <= 12'h0;
    end
    copyEnabledReg <= preDisplayArea & _T_365;
    _T_373 <= backMemoryRestoreCounter[10:0];
    _T_375 <= io_backBufferWriteAddress;
    _T_378 <= backMemoryRestoreCounter < 12'h800;
    _T_379 <= io_backBufferWriteEnable;
    _T_382 <= io_backBufferWriteData;
    _T_385 <= backMemoryCopyCounter[10:0];
    _T_393 <= backMemoryRestoreCounter[10:0];
    _T_395 <= io_backBufferWriteAddress;
    _T_398 <= backMemoryRestoreCounter < 12'h800;
    _T_399 <= io_backBufferWriteEnable;
    _T_402 <= io_backBufferWriteData;
    _T_405 <= backMemoryCopyCounter[10:0];
    _T_412 <= backBufferMemories_0_io_dataRead;
    _T_415 <= backBufferMemories_1_io_dataRead;
    if (fullBackgroundColor_0[6]) begin
      if (fullBackgroundColor_1[6]) begin
        pixelColorBack <= 6'h0;
      end else begin
        pixelColorBack <= fullBackgroundColor_1[5:0];
      end
    end else begin
      pixelColorBack <= fullBackgroundColor_0[5:0];
    end
    _T_3497 <= spriteMemories_0_io_dataRead[5:0];
    _T_3498_0 <= _T_3498_1;
    _T_3498_1 <= spriteVisibleReg_0;
    _T_3499_0 <= _T_3499_1;
    _T_3499_1 <= _T_440 & _T_441;
    _T_3502 <= spriteMemories_0_io_dataRead[6];
    _T_3506 <= spriteMemories_1_io_dataRead[5:0];
    _T_3507_0 <= _T_3507_1;
    _T_3507_1 <= spriteVisibleReg_1;
    _T_3508_0 <= _T_3508_1;
    _T_3508_1 <= _T_459 & _T_460;
    _T_3511 <= spriteMemories_1_io_dataRead[6];
    _T_3515 <= spriteMemories_2_io_dataRead[5:0];
    _T_3516_0 <= _T_3516_1;
    _T_3516_1 <= spriteVisibleReg_2;
    _T_3517_0 <= _T_3517_1;
    _T_3517_1 <= _T_478 & _T_479;
    _T_3520 <= spriteMemories_2_io_dataRead[6];
    _T_3524 <= spriteMemories_3_io_dataRead[5:0];
    _T_3525_0 <= _T_3525_1;
    _T_3525_1 <= spriteVisibleReg_3;
    _T_3526_0 <= _T_3526_1;
    _T_3526_1 <= _T_497 & _T_498;
    _T_3529 <= spriteMemories_3_io_dataRead[6];
    _T_3533 <= spriteMemories_4_io_dataRead[5:0];
    _T_3534_0 <= _T_3534_1;
    _T_3534_1 <= spriteVisibleReg_4;
    _T_3535_0 <= _T_3535_1;
    _T_3535_1 <= _T_516 & _T_517;
    _T_3538 <= spriteMemories_4_io_dataRead[6];
    _T_3542 <= spriteMemories_5_io_dataRead[5:0];
    _T_3543_0 <= _T_3543_1;
    _T_3543_1 <= spriteVisibleReg_5;
    _T_3544_0 <= _T_3544_1;
    _T_3544_1 <= _T_535 & _T_536;
    _T_3547 <= spriteMemories_5_io_dataRead[6];
    _T_3551 <= spriteMemories_6_io_dataRead[5:0];
    _T_3552_0 <= _T_3552_1;
    _T_3552_1 <= spriteVisibleReg_6;
    _T_3553_0 <= _T_3553_1;
    _T_3553_1 <= _T_554 & _T_555;
    _T_3556 <= spriteMemories_6_io_dataRead[6];
    _T_3560 <= spriteMemories_7_io_dataRead[5:0];
    _T_3561_0 <= _T_3561_1;
    _T_3561_1 <= spriteVisibleReg_7;
    _T_3562_0 <= _T_3562_1;
    _T_3562_1 <= _T_573 & _T_574;
    _T_3565 <= spriteMemories_7_io_dataRead[6];
    _T_3569 <= spriteMemories_8_io_dataRead[5:0];
    _T_3570_0 <= _T_3570_1;
    _T_3570_1 <= spriteVisibleReg_8;
    _T_3571_0 <= _T_3571_1;
    _T_3571_1 <= _T_592 & _T_593;
    _T_3574 <= spriteMemories_8_io_dataRead[6];
    _T_3578 <= spriteMemories_9_io_dataRead[5:0];
    _T_3579_0 <= _T_3579_1;
    _T_3579_1 <= spriteVisibleReg_9;
    _T_3580_0 <= _T_3580_1;
    _T_3580_1 <= _T_611 & _T_612;
    _T_3583 <= spriteMemories_9_io_dataRead[6];
    _T_3587 <= spriteMemories_10_io_dataRead[5:0];
    _T_3588_0 <= _T_3588_1;
    _T_3588_1 <= spriteVisibleReg_10;
    _T_3589_0 <= _T_3589_1;
    _T_3589_1 <= _T_630 & _T_631;
    _T_3592 <= spriteMemories_10_io_dataRead[6];
    _T_3596 <= spriteMemories_11_io_dataRead[5:0];
    _T_3597_0 <= _T_3597_1;
    _T_3597_1 <= spriteVisibleReg_11;
    _T_3598_0 <= _T_3598_1;
    _T_3598_1 <= _T_649 & _T_650;
    _T_3601 <= spriteMemories_11_io_dataRead[6];
    _T_3605 <= spriteMemories_12_io_dataRead[5:0];
    _T_3606_0 <= _T_3606_1;
    _T_3606_1 <= spriteVisibleReg_12;
    _T_3607_0 <= _T_3607_1;
    _T_3607_1 <= _T_668 & _T_669;
    _T_3610 <= spriteMemories_12_io_dataRead[6];
    _T_3614 <= spriteMemories_13_io_dataRead[5:0];
    _T_3615_0 <= _T_3615_1;
    _T_3615_1 <= spriteVisibleReg_13;
    _T_3616_0 <= _T_3616_1;
    _T_3616_1 <= _T_687 & _T_688;
    _T_3619 <= spriteMemories_13_io_dataRead[6];
    _T_3623 <= spriteMemories_14_io_dataRead[5:0];
    _T_3624_0 <= _T_3624_1;
    _T_3624_1 <= spriteVisibleReg_14;
    _T_3625_0 <= _T_3625_1;
    _T_3625_1 <= _T_706 & _T_707;
    _T_3628 <= spriteMemories_14_io_dataRead[6];
    _T_3632 <= spriteMemories_15_io_dataRead[5:0];
    _T_3633_0 <= _T_3633_1;
    _T_3633_1 <= spriteVisibleReg_15;
    _T_3634_0 <= _T_3634_1;
    _T_3634_1 <= _T_725 & _T_726;
    _T_3637 <= spriteMemories_15_io_dataRead[6];
    _T_3641 <= spriteMemories_16_io_dataRead[5:0];
    _T_3642_0 <= _T_3642_1;
    _T_3642_1 <= spriteVisibleReg_16;
    _T_3643_0 <= _T_3643_1;
    _T_3643_1 <= _T_744 & _T_745;
    _T_3646 <= spriteMemories_16_io_dataRead[6];
    _T_3650 <= spriteMemories_17_io_dataRead[5:0];
    _T_3651_0 <= _T_3651_1;
    _T_3651_1 <= spriteVisibleReg_17;
    _T_3652_0 <= _T_3652_1;
    _T_3652_1 <= _T_763 & _T_764;
    _T_3655 <= spriteMemories_17_io_dataRead[6];
    _T_3659 <= spriteMemories_18_io_dataRead[5:0];
    _T_3660_0 <= _T_3660_1;
    _T_3660_1 <= spriteVisibleReg_18;
    _T_3661_0 <= _T_3661_1;
    _T_3661_1 <= _T_782 & _T_783;
    _T_3664 <= spriteMemories_18_io_dataRead[6];
    _T_3668 <= spriteMemories_19_io_dataRead[5:0];
    _T_3669_0 <= _T_3669_1;
    _T_3669_1 <= spriteVisibleReg_19;
    _T_3670_0 <= _T_3670_1;
    _T_3670_1 <= _T_801 & _T_802;
    _T_3673 <= spriteMemories_19_io_dataRead[6];
    _T_3677 <= spriteMemories_20_io_dataRead[5:0];
    _T_3678_0 <= _T_3678_1;
    _T_3678_1 <= spriteVisibleReg_20;
    _T_3679_0 <= _T_3679_1;
    _T_3679_1 <= _T_820 & _T_821;
    _T_3682 <= spriteMemories_20_io_dataRead[6];
    _T_3686 <= spriteMemories_21_io_dataRead[5:0];
    _T_3687_0 <= _T_3687_1;
    _T_3687_1 <= spriteVisibleReg_21;
    _T_3688_0 <= _T_3688_1;
    _T_3688_1 <= _T_839 & _T_840;
    _T_3691 <= spriteMemories_21_io_dataRead[6];
    _T_3695 <= spriteMemories_22_io_dataRead[5:0];
    _T_3696_0 <= _T_3696_1;
    _T_3696_1 <= spriteVisibleReg_22;
    _T_3697_0 <= _T_3697_1;
    _T_3697_1 <= _T_858 & _T_859;
    _T_3700 <= spriteMemories_22_io_dataRead[6];
    _T_3704 <= spriteMemories_23_io_dataRead[5:0];
    _T_3705_0 <= _T_3705_1;
    _T_3705_1 <= spriteVisibleReg_23;
    _T_3706_0 <= _T_3706_1;
    _T_3706_1 <= _T_877 & _T_878;
    _T_3709 <= spriteMemories_23_io_dataRead[6];
    _T_3713 <= spriteMemories_24_io_dataRead[5:0];
    _T_3714_0 <= _T_3714_1;
    _T_3714_1 <= spriteVisibleReg_24;
    _T_3715_0 <= _T_3715_1;
    _T_3715_1 <= _T_896 & _T_897;
    _T_3718 <= spriteMemories_24_io_dataRead[6];
    _T_3722 <= spriteMemories_25_io_dataRead[5:0];
    _T_3723_0 <= _T_3723_1;
    _T_3723_1 <= spriteVisibleReg_25;
    _T_3724_0 <= _T_3724_1;
    _T_3724_1 <= _T_915 & _T_916;
    _T_3727 <= spriteMemories_25_io_dataRead[6];
    _T_3731 <= spriteMemories_26_io_dataRead[5:0];
    _T_3732_0 <= _T_3732_1;
    _T_3732_1 <= spriteVisibleReg_26;
    _T_3733_0 <= _T_3733_1;
    _T_3733_1 <= _T_934 & _T_935;
    _T_3736 <= spriteMemories_26_io_dataRead[6];
    _T_3740 <= spriteMemories_27_io_dataRead[5:0];
    _T_3741_0 <= _T_3741_1;
    _T_3741_1 <= spriteVisibleReg_27;
    _T_3742_0 <= _T_3742_1;
    _T_3742_1 <= _T_953 & _T_954;
    _T_3745 <= spriteMemories_27_io_dataRead[6];
    _T_3749 <= spriteMemories_28_io_dataRead[5:0];
    _T_3750_0 <= _T_3750_1;
    _T_3750_1 <= spriteVisibleReg_28;
    _T_3751_0 <= _T_3751_1;
    _T_3751_1 <= _T_972 & _T_973;
    _T_3754 <= spriteMemories_28_io_dataRead[6];
    _T_3758 <= spriteMemories_29_io_dataRead[5:0];
    _T_3759_0 <= _T_3759_1;
    _T_3759_1 <= spriteVisibleReg_29;
    _T_3760_0 <= _T_3760_1;
    _T_3760_1 <= _T_991 & _T_992;
    _T_3763 <= spriteMemories_29_io_dataRead[6];
    _T_3767 <= spriteMemories_30_io_dataRead[5:0];
    _T_3768_0 <= _T_3768_1;
    _T_3768_1 <= spriteVisibleReg_30;
    _T_3769_0 <= _T_3769_1;
    _T_3769_1 <= _T_1010 & _T_1011;
    _T_3772 <= spriteMemories_30_io_dataRead[6];
    _T_3776 <= spriteMemories_31_io_dataRead[5:0];
    _T_3777_0 <= _T_3777_1;
    _T_3777_1 <= spriteVisibleReg_31;
    _T_3778_0 <= _T_3778_1;
    _T_3778_1 <= _T_1029 & _T_1030;
    _T_3781 <= spriteMemories_31_io_dataRead[6];
    _T_3785 <= spriteMemories_32_io_dataRead[5:0];
    _T_3786_0 <= _T_3786_1;
    _T_3786_1 <= spriteVisibleReg_32;
    _T_3787_0 <= _T_3787_1;
    _T_3787_1 <= _T_1048 & _T_1049;
    _T_3790 <= spriteMemories_32_io_dataRead[6];
    _T_3794 <= spriteMemories_33_io_dataRead[5:0];
    _T_3795_0 <= _T_3795_1;
    _T_3795_1 <= spriteVisibleReg_33;
    _T_3796_0 <= _T_3796_1;
    _T_3796_1 <= _T_1067 & _T_1068;
    _T_3799 <= spriteMemories_33_io_dataRead[6];
    _T_3803 <= spriteMemories_34_io_dataRead[5:0];
    _T_3805_0 <= _T_3805_1;
    _T_3805_1 <= _T_1086 & _T_1087;
    _T_3808 <= spriteMemories_34_io_dataRead[6];
    _T_3812 <= spriteMemories_35_io_dataRead[5:0];
    _T_3814_0 <= _T_3814_1;
    _T_3814_1 <= _T_1105 & _T_1106;
    _T_3817 <= spriteMemories_35_io_dataRead[6];
    _T_3821 <= spriteMemories_36_io_dataRead[5:0];
    _T_3823_0 <= _T_3823_1;
    _T_3823_1 <= _T_1124 & _T_1125;
    _T_3826 <= spriteMemories_36_io_dataRead[6];
    _T_3830 <= spriteMemories_37_io_dataRead[5:0];
    _T_3832_0 <= _T_3832_1;
    _T_3832_1 <= _T_1143 & _T_1144;
    _T_3835 <= spriteMemories_37_io_dataRead[6];
    _T_3839 <= spriteMemories_38_io_dataRead[5:0];
    _T_3841_0 <= _T_3841_1;
    _T_3841_1 <= _T_1162 & _T_1163;
    _T_3844 <= spriteMemories_38_io_dataRead[6];
    _T_3848 <= spriteMemories_39_io_dataRead[5:0];
    _T_3850_0 <= _T_3850_1;
    _T_3850_1 <= _T_1181 & _T_1182;
    _T_3853 <= spriteMemories_39_io_dataRead[6];
    _T_3857 <= spriteMemories_40_io_dataRead[5:0];
    _T_3859_0 <= _T_3859_1;
    _T_3859_1 <= _T_1200 & _T_1201;
    _T_3862 <= spriteMemories_40_io_dataRead[6];
    _T_3866 <= spriteMemories_41_io_dataRead[5:0];
    _T_3867_0 <= _T_3867_1;
    _T_3867_1 <= spriteVisibleReg_41;
    _T_3868_0 <= _T_3868_1;
    _T_3868_1 <= _T_1219 & _T_1220;
    _T_3871 <= spriteMemories_41_io_dataRead[6];
    _T_3875 <= spriteMemories_42_io_dataRead[5:0];
    _T_3876_0 <= _T_3876_1;
    _T_3876_1 <= spriteVisibleReg_42;
    _T_3877_0 <= _T_3877_1;
    _T_3877_1 <= _T_1238 & _T_1239;
    _T_3880 <= spriteMemories_42_io_dataRead[6];
    _T_3884 <= spriteMemories_43_io_dataRead[5:0];
    _T_3885_0 <= _T_3885_1;
    _T_3885_1 <= spriteVisibleReg_43;
    _T_3886_0 <= _T_3886_1;
    _T_3886_1 <= _T_1257 & _T_1258;
    _T_3889 <= spriteMemories_43_io_dataRead[6];
    _T_3893 <= spriteMemories_44_io_dataRead[5:0];
    _T_3894_0 <= _T_3894_1;
    _T_3894_1 <= spriteVisibleReg_44;
    _T_3895_0 <= _T_3895_1;
    _T_3895_1 <= _T_1276 & _T_1277;
    _T_3898 <= spriteMemories_44_io_dataRead[6];
    _T_3902 <= spriteMemories_45_io_dataRead[5:0];
    _T_3903_0 <= _T_3903_1;
    _T_3903_1 <= spriteVisibleReg_45;
    _T_3904_0 <= _T_3904_1;
    _T_3904_1 <= _T_1295 & _T_1296;
    _T_3907 <= spriteMemories_45_io_dataRead[6];
    _T_3911 <= spriteMemories_46_io_dataRead[5:0];
    _T_3912_0 <= _T_3912_1;
    _T_3912_1 <= spriteVisibleReg_46;
    _T_3913_0 <= _T_3913_1;
    _T_3913_1 <= _T_1314 & _T_1315;
    _T_3916 <= spriteMemories_46_io_dataRead[6];
    _T_3920 <= spriteMemories_47_io_dataRead[5:0];
    _T_3921_0 <= _T_3921_1;
    _T_3921_1 <= spriteVisibleReg_47;
    _T_3922_0 <= _T_3922_1;
    _T_3922_1 <= _T_1333 & _T_1334;
    _T_3925 <= spriteMemories_47_io_dataRead[6];
    _T_3929 <= spriteMemories_48_io_dataRead[5:0];
    _T_3930_0 <= _T_3930_1;
    _T_3930_1 <= spriteVisibleReg_48;
    _T_3931_0 <= _T_3931_1;
    _T_3931_1 <= _T_1352 & _T_1353;
    _T_3934 <= spriteMemories_48_io_dataRead[6];
    _T_3938 <= spriteMemories_49_io_dataRead[5:0];
    _T_3939_0 <= _T_3939_1;
    _T_3939_1 <= spriteVisibleReg_49;
    _T_3940_0 <= _T_3940_1;
    _T_3940_1 <= _T_1371 & _T_1372;
    _T_3943 <= spriteMemories_49_io_dataRead[6];
    _T_3947 <= spriteMemories_50_io_dataRead[5:0];
    _T_3948_0 <= _T_3948_1;
    _T_3948_1 <= spriteVisibleReg_50;
    _T_3949_0 <= _T_3949_1;
    _T_3949_1 <= _T_1390 & _T_1391;
    _T_3952 <= spriteMemories_50_io_dataRead[6];
    _T_3956 <= spriteMemories_51_io_dataRead[5:0];
    _T_3957_0 <= _T_3957_1;
    _T_3957_1 <= spriteVisibleReg_51;
    _T_3958_0 <= _T_3958_1;
    _T_3958_1 <= _T_1409 & _T_1410;
    _T_3961 <= spriteMemories_51_io_dataRead[6];
    _T_3965 <= spriteMemories_52_io_dataRead[5:0];
    _T_3967_0 <= _T_3967_1;
    _T_3967_1 <= _T_1428 & _T_1429;
    _T_3970 <= spriteMemories_52_io_dataRead[6];
    _T_3974 <= spriteMemories_53_io_dataRead[5:0];
    _T_3976_0 <= _T_3976_1;
    _T_3976_1 <= _T_1447 & _T_1448;
    _T_3979 <= spriteMemories_53_io_dataRead[6];
    _T_3983 <= spriteMemories_54_io_dataRead[5:0];
    _T_3985_0 <= _T_3985_1;
    _T_3985_1 <= _T_1466 & _T_1467;
    _T_3988 <= spriteMemories_54_io_dataRead[6];
    _T_3992 <= spriteMemories_55_io_dataRead[5:0];
    _T_3993_0 <= _T_3993_1;
    _T_3993_1 <= spriteVisibleReg_55;
    _T_3994_0 <= _T_3994_1;
    _T_3994_1 <= _T_1485 & _T_1486;
    _T_3997 <= spriteMemories_55_io_dataRead[6];
    _T_4001 <= spriteMemories_56_io_dataRead[5:0];
    _T_4002_0 <= _T_4002_1;
    _T_4002_1 <= spriteVisibleReg_56;
    _T_4003_0 <= _T_4003_1;
    _T_4003_1 <= _T_1504 & _T_1505;
    _T_4006 <= spriteMemories_56_io_dataRead[6];
    _T_4010 <= spriteMemories_57_io_dataRead[5:0];
    _T_4011_0 <= _T_4011_1;
    _T_4011_1 <= spriteVisibleReg_57;
    _T_4012_0 <= _T_4012_1;
    _T_4012_1 <= _T_1523 & _T_1524;
    _T_4015 <= spriteMemories_57_io_dataRead[6];
    _T_4019 <= spriteMemories_58_io_dataRead[5:0];
    _T_4021_0 <= _T_4021_1;
    _T_4021_1 <= _T_1542 & _T_1543;
    _T_4024 <= spriteMemories_58_io_dataRead[6];
    _T_4028 <= spriteMemories_59_io_dataRead[5:0];
    _T_4030_0 <= _T_4030_1;
    _T_4030_1 <= _T_1561 & _T_1562;
    _T_4033 <= spriteMemories_59_io_dataRead[6];
    _T_4037 <= spriteMemories_60_io_dataRead[5:0];
    _T_4039_0 <= _T_4039_1;
    _T_4039_1 <= _T_1580 & _T_1581;
    _T_4042 <= spriteMemories_60_io_dataRead[6];
    _T_4046 <= spriteMemories_61_io_dataRead[5:0];
    _T_4047_0 <= _T_4047_1;
    _T_4047_1 <= spriteVisibleReg_61;
    _T_4048_0 <= _T_4048_1;
    _T_4048_1 <= _T_1599 & _T_1600;
    _T_4051 <= spriteMemories_61_io_dataRead[6];
    _T_4055 <= spriteMemories_62_io_dataRead[5:0];
    _T_4056_0 <= _T_4056_1;
    _T_4056_1 <= spriteVisibleReg_62;
    _T_4057_0 <= _T_4057_1;
    _T_4057_1 <= _T_1618 & _T_1619;
    _T_4060 <= spriteMemories_62_io_dataRead[6];
    _T_4064 <= spriteMemories_63_io_dataRead[5:0];
    _T_4065_0 <= _T_4065_1;
    _T_4065_1 <= spriteVisibleReg_63;
    _T_4066_0 <= _T_4066_1;
    _T_4066_1 <= _T_1637 & _T_1638;
    _T_4069 <= spriteMemories_63_io_dataRead[6];
    _T_4073 <= spriteMemories_64_io_dataRead[5:0];
    _T_4074_0 <= _T_4074_1;
    _T_4074_1 <= spriteVisibleReg_64;
    _T_4075_0 <= _T_4075_1;
    _T_4075_1 <= _T_1656 & _T_1657;
    _T_4078 <= spriteMemories_64_io_dataRead[6];
    _T_4082 <= spriteMemories_65_io_dataRead[5:0];
    _T_4083_0 <= _T_4083_1;
    _T_4083_1 <= spriteVisibleReg_65;
    _T_4084_0 <= _T_4084_1;
    _T_4084_1 <= _T_1675 & _T_1657;
    _T_4087 <= spriteMemories_65_io_dataRead[6];
    _T_4091 <= spriteMemories_66_io_dataRead[5:0];
    _T_4092_0 <= _T_4092_1;
    _T_4092_1 <= spriteVisibleReg_66;
    _T_4093_0 <= _T_4093_1;
    _T_4093_1 <= _T_1694 & _T_1657;
    _T_4096 <= spriteMemories_66_io_dataRead[6];
    _T_4100 <= spriteMemories_67_io_dataRead[5:0];
    _T_4102_0 <= _T_4102_1;
    _T_4102_1 <= _T_1713 & _T_1657;
    _T_4105 <= spriteMemories_67_io_dataRead[6];
    _T_4109 <= spriteMemories_68_io_dataRead[5:0];
    _T_4111_0 <= _T_4111_1;
    _T_4111_1 <= _T_1732 & _T_1657;
    _T_4114 <= spriteMemories_68_io_dataRead[6];
    _T_4118 <= spriteMemories_69_io_dataRead[5:0];
    _T_4120_0 <= _T_4120_1;
    _T_4120_1 <= _T_1751 & _T_1657;
    _T_4123 <= spriteMemories_69_io_dataRead[6];
    _T_4127 <= spriteMemories_70_io_dataRead[5:0];
    _T_4128_0 <= _T_4128_1;
    _T_4128_1 <= spriteVisibleReg_70;
    _T_4129_0 <= _T_4129_1;
    _T_4129_1 <= _T_1770 & _T_1771;
    _T_4132 <= spriteMemories_70_io_dataRead[6];
    _T_4136 <= spriteMemories_71_io_dataRead[5:0];
    _T_4137_0 <= _T_4137_1;
    _T_4137_1 <= spriteVisibleReg_71;
    _T_4138_0 <= _T_4138_1;
    _T_4138_1 <= _T_1789 & _T_1790;
    _T_4141 <= spriteMemories_71_io_dataRead[6];
    _T_4145 <= spriteMemories_72_io_dataRead[5:0];
    _T_4146_0 <= _T_4146_1;
    _T_4146_1 <= spriteVisibleReg_72;
    _T_4147_0 <= _T_4147_1;
    _T_4147_1 <= _T_1808 & _T_1809;
    _T_4150 <= spriteMemories_72_io_dataRead[6];
    _T_4154 <= spriteMemories_73_io_dataRead[5:0];
    _T_4156_0 <= _T_4156_1;
    _T_4156_1 <= _T_1827 & _T_1828;
    _T_4159 <= spriteMemories_73_io_dataRead[6];
    _T_4163 <= spriteMemories_74_io_dataRead[5:0];
    _T_4165_0 <= _T_4165_1;
    _T_4165_1 <= _T_1846 & _T_1847;
    _T_4168 <= spriteMemories_74_io_dataRead[6];
    _T_4172 <= spriteMemories_75_io_dataRead[5:0];
    _T_4174_0 <= _T_4174_1;
    _T_4174_1 <= _T_1865 & _T_1866;
    _T_4177 <= spriteMemories_75_io_dataRead[6];
    _T_4181 <= spriteMemories_76_io_dataRead[5:0];
    _T_4183_0 <= _T_4183_1;
    _T_4183_1 <= _T_1884 & _T_1885;
    _T_4186 <= spriteMemories_76_io_dataRead[6];
    _T_4190 <= spriteMemories_77_io_dataRead[5:0];
    _T_4192_0 <= _T_4192_1;
    _T_4192_1 <= _T_1903 & _T_1904;
    _T_4195 <= spriteMemories_77_io_dataRead[6];
    _T_4199 <= spriteMemories_78_io_dataRead[5:0];
    _T_4201_0 <= _T_4201_1;
    _T_4201_1 <= _T_1922 & _T_1923;
    _T_4204 <= spriteMemories_78_io_dataRead[6];
    _T_4208 <= spriteMemories_79_io_dataRead[5:0];
    _T_4210_0 <= _T_4210_1;
    _T_4210_1 <= _T_1941 & _T_1942;
    _T_4213 <= spriteMemories_79_io_dataRead[6];
    _T_4217 <= spriteMemories_80_io_dataRead[5:0];
    _T_4219_0 <= _T_4219_1;
    _T_4219_1 <= _T_1960 & _T_1961;
    _T_4222 <= spriteMemories_80_io_dataRead[6];
    _T_4226 <= spriteMemories_81_io_dataRead[5:0];
    _T_4228_0 <= _T_4228_1;
    _T_4228_1 <= _T_1979 & _T_1980;
    _T_4231 <= spriteMemories_81_io_dataRead[6];
    _T_4235 <= spriteMemories_82_io_dataRead[5:0];
    _T_4237_0 <= _T_4237_1;
    _T_4237_1 <= _T_1998 & _T_1999;
    _T_4240 <= spriteMemories_82_io_dataRead[6];
    _T_4244 <= spriteMemories_83_io_dataRead[5:0];
    _T_4246_0 <= _T_4246_1;
    _T_4246_1 <= _T_2017 & _T_2018;
    _T_4249 <= spriteMemories_83_io_dataRead[6];
    _T_4253 <= spriteMemories_84_io_dataRead[5:0];
    _T_4255_0 <= _T_4255_1;
    _T_4255_1 <= _T_2036 & _T_2037;
    _T_4258 <= spriteMemories_84_io_dataRead[6];
    _T_4262 <= spriteMemories_85_io_dataRead[5:0];
    _T_4264_0 <= _T_4264_1;
    _T_4264_1 <= _T_2055 & _T_2056;
    _T_4267 <= spriteMemories_85_io_dataRead[6];
    _T_4271 <= spriteMemories_86_io_dataRead[5:0];
    _T_4273_0 <= _T_4273_1;
    _T_4273_1 <= _T_2074 & _T_2075;
    _T_4276 <= spriteMemories_86_io_dataRead[6];
    _T_4280 <= spriteMemories_87_io_dataRead[5:0];
    _T_4282_0 <= _T_4282_1;
    _T_4282_1 <= _T_2093 & _T_2094;
    _T_4285 <= spriteMemories_87_io_dataRead[6];
    _T_4289 <= spriteMemories_88_io_dataRead[5:0];
    _T_4291_0 <= _T_4291_1;
    _T_4291_1 <= _T_2112 & _T_2113;
    _T_4294 <= spriteMemories_88_io_dataRead[6];
    _T_4298 <= spriteMemories_89_io_dataRead[5:0];
    _T_4300_0 <= _T_4300_1;
    _T_4300_1 <= _T_2131 & _T_2132;
    _T_4303 <= spriteMemories_89_io_dataRead[6];
    _T_4307 <= spriteMemories_90_io_dataRead[5:0];
    _T_4309_0 <= _T_4309_1;
    _T_4309_1 <= _T_2150 & _T_2151;
    _T_4312 <= spriteMemories_90_io_dataRead[6];
    _T_4316 <= spriteMemories_91_io_dataRead[5:0];
    _T_4318_0 <= _T_4318_1;
    _T_4318_1 <= _T_2169 & _T_2170;
    _T_4321 <= spriteMemories_91_io_dataRead[6];
    _T_4325 <= spriteMemories_92_io_dataRead[5:0];
    _T_4327_0 <= _T_4327_1;
    _T_4327_1 <= _T_2188 & _T_2189;
    _T_4330 <= spriteMemories_92_io_dataRead[6];
    _T_4334 <= spriteMemories_93_io_dataRead[5:0];
    _T_4336_0 <= _T_4336_1;
    _T_4336_1 <= _T_2207 & _T_2208;
    _T_4339 <= spriteMemories_93_io_dataRead[6];
    _T_4343 <= spriteMemories_94_io_dataRead[5:0];
    _T_4345_0 <= _T_4345_1;
    _T_4345_1 <= _T_2226 & _T_2227;
    _T_4348 <= spriteMemories_94_io_dataRead[6];
    _T_4352 <= spriteMemories_95_io_dataRead[5:0];
    _T_4354_0 <= _T_4354_1;
    _T_4354_1 <= _T_2245 & _T_2246;
    _T_4357 <= spriteMemories_95_io_dataRead[6];
    _T_4361 <= spriteMemories_96_io_dataRead[5:0];
    _T_4363_0 <= _T_4363_1;
    _T_4363_1 <= _T_2264 & _T_2265;
    _T_4366 <= spriteMemories_96_io_dataRead[6];
    _T_4370 <= spriteMemories_97_io_dataRead[5:0];
    _T_4372_0 <= _T_4372_1;
    _T_4372_1 <= _T_2283 & _T_2284;
    _T_4375 <= spriteMemories_97_io_dataRead[6];
    _T_4379 <= spriteMemories_98_io_dataRead[5:0];
    _T_4381_0 <= _T_4381_1;
    _T_4381_1 <= _T_2302 & _T_2303;
    _T_4384 <= spriteMemories_98_io_dataRead[6];
    _T_4388 <= spriteMemories_99_io_dataRead[5:0];
    _T_4390_0 <= _T_4390_1;
    _T_4390_1 <= _T_2321 & _T_2322;
    _T_4393 <= spriteMemories_99_io_dataRead[6];
    _T_4397 <= spriteMemories_100_io_dataRead[5:0];
    _T_4399_0 <= _T_4399_1;
    _T_4399_1 <= _T_2340 & _T_2341;
    _T_4402 <= spriteMemories_100_io_dataRead[6];
    _T_4406 <= spriteMemories_101_io_dataRead[5:0];
    _T_4408_0 <= _T_4408_1;
    _T_4408_1 <= _T_2359 & _T_2360;
    _T_4411 <= spriteMemories_101_io_dataRead[6];
    _T_4415 <= spriteMemories_102_io_dataRead[5:0];
    _T_4417_0 <= _T_4417_1;
    _T_4417_1 <= _T_2378 & _T_2379;
    _T_4420 <= spriteMemories_102_io_dataRead[6];
    _T_4424 <= spriteMemories_103_io_dataRead[5:0];
    _T_4426_0 <= _T_4426_1;
    _T_4426_1 <= _T_2397 & _T_2398;
    _T_4429 <= spriteMemories_103_io_dataRead[6];
    _T_4433 <= spriteMemories_104_io_dataRead[5:0];
    _T_4435_0 <= _T_4435_1;
    _T_4435_1 <= _T_2416 & _T_2417;
    _T_4438 <= spriteMemories_104_io_dataRead[6];
    _T_4442 <= spriteMemories_105_io_dataRead[5:0];
    _T_4444_0 <= _T_4444_1;
    _T_4444_1 <= _T_2435 & _T_2436;
    _T_4447 <= spriteMemories_105_io_dataRead[6];
    _T_4451 <= spriteMemories_106_io_dataRead[5:0];
    _T_4453_0 <= _T_4453_1;
    _T_4453_1 <= _T_2454 & _T_2455;
    _T_4456 <= spriteMemories_106_io_dataRead[6];
    _T_4460 <= spriteMemories_107_io_dataRead[5:0];
    _T_4462_0 <= _T_4462_1;
    _T_4462_1 <= _T_2473 & _T_2474;
    _T_4465 <= spriteMemories_107_io_dataRead[6];
    _T_4469 <= spriteMemories_108_io_dataRead[5:0];
    _T_4471_0 <= _T_4471_1;
    _T_4471_1 <= _T_2492 & _T_2493;
    _T_4474 <= spriteMemories_108_io_dataRead[6];
    _T_4478 <= spriteMemories_109_io_dataRead[5:0];
    _T_4480_0 <= _T_4480_1;
    _T_4480_1 <= _T_2511 & _T_2512;
    _T_4483 <= spriteMemories_109_io_dataRead[6];
    _T_4487 <= spriteMemories_110_io_dataRead[5:0];
    _T_4489_0 <= _T_4489_1;
    _T_4489_1 <= _T_2530 & _T_2531;
    _T_4492 <= spriteMemories_110_io_dataRead[6];
    _T_4496 <= spriteMemories_111_io_dataRead[5:0];
    _T_4498_0 <= _T_4498_1;
    _T_4498_1 <= _T_2549 & _T_2550;
    _T_4501 <= spriteMemories_111_io_dataRead[6];
    _T_4505 <= spriteMemories_112_io_dataRead[5:0];
    _T_4507_0 <= _T_4507_1;
    _T_4507_1 <= _T_2568 & _T_2569;
    _T_4510 <= spriteMemories_112_io_dataRead[6];
    _T_4514 <= spriteMemories_113_io_dataRead[5:0];
    _T_4516_0 <= _T_4516_1;
    _T_4516_1 <= _T_2587 & _T_2588;
    _T_4519 <= spriteMemories_113_io_dataRead[6];
    _T_4523 <= spriteMemories_114_io_dataRead[5:0];
    _T_4525_0 <= _T_4525_1;
    _T_4525_1 <= _T_2606 & _T_2607;
    _T_4528 <= spriteMemories_114_io_dataRead[6];
    _T_4532 <= spriteMemories_115_io_dataRead[5:0];
    _T_4534_0 <= _T_4534_1;
    _T_4534_1 <= _T_2625 & _T_2626;
    _T_4537 <= spriteMemories_115_io_dataRead[6];
    _T_4541 <= spriteMemories_116_io_dataRead[5:0];
    _T_4543_0 <= _T_4543_1;
    _T_4543_1 <= _T_2644 & _T_2645;
    _T_4546 <= spriteMemories_116_io_dataRead[6];
    _T_4550 <= spriteMemories_117_io_dataRead[5:0];
    _T_4552_0 <= _T_4552_1;
    _T_4552_1 <= _T_2663 & _T_2664;
    _T_4555 <= spriteMemories_117_io_dataRead[6];
    _T_4559 <= spriteMemories_118_io_dataRead[5:0];
    _T_4561_0 <= _T_4561_1;
    _T_4561_1 <= _T_2682 & _T_2683;
    _T_4564 <= spriteMemories_118_io_dataRead[6];
    _T_4568 <= spriteMemories_119_io_dataRead[5:0];
    _T_4570_0 <= _T_4570_1;
    _T_4570_1 <= _T_2701 & _T_2702;
    _T_4573 <= spriteMemories_119_io_dataRead[6];
    _T_4577 <= spriteMemories_120_io_dataRead[5:0];
    _T_4579_0 <= _T_4579_1;
    _T_4579_1 <= _T_2720 & _T_2721;
    _T_4582 <= spriteMemories_120_io_dataRead[6];
    _T_4586 <= spriteMemories_121_io_dataRead[5:0];
    _T_4588_0 <= _T_4588_1;
    _T_4588_1 <= _T_2739 & _T_2740;
    _T_4591 <= spriteMemories_121_io_dataRead[6];
    _T_4595 <= spriteMemories_122_io_dataRead[5:0];
    _T_4597_0 <= _T_4597_1;
    _T_4597_1 <= _T_2758 & _T_2759;
    _T_4600 <= spriteMemories_122_io_dataRead[6];
    _T_4604 <= spriteMemories_123_io_dataRead[5:0];
    _T_4606_0 <= _T_4606_1;
    _T_4606_1 <= _T_2777 & _T_2778;
    _T_4609 <= spriteMemories_123_io_dataRead[6];
    _T_4613 <= spriteMemories_124_io_dataRead[5:0];
    _T_4615_0 <= _T_4615_1;
    _T_4615_1 <= _T_2796 & _T_2797;
    _T_4618 <= spriteMemories_124_io_dataRead[6];
    _T_4622 <= spriteMemories_125_io_dataRead[5:0];
    _T_4624_0 <= _T_4624_1;
    _T_4624_1 <= _T_2815 & _T_2816;
    _T_4627 <= spriteMemories_125_io_dataRead[6];
    _T_4631 <= spriteMemories_126_io_dataRead[5:0];
    _T_4633_0 <= _T_4633_1;
    _T_4633_1 <= _T_2834 & _T_2835;
    _T_4636 <= spriteMemories_126_io_dataRead[6];
    _T_4640 <= spriteMemories_127_io_dataRead[5:0];
    _T_4642_0 <= _T_4642_1;
    _T_4642_1 <= _T_2853 & _T_2854;
    _T_4645 <= spriteMemories_127_io_dataRead[6];
    pixelColorSprite <= multiHotPriortyReductionTree_io_dataOutput;
    pixelColorSpriteValid <= multiHotPriortyReductionTree_io_selectOutput;
    _T_4648_0 <= _T_4648_1;
    _T_4648_1 <= _T_4648_2;
    _T_4648_2 <= _T_17 & _T_18;
    _T_4655 <= {pixelColourVGA[5:4],pixelColourVGA[5:4]};
    _T_4656 <= {pixelColourVGA[3:2],pixelColourVGA[3:2]};
    _T_4657 <= {pixelColourVGA[1:0],pixelColourVGA[1:0]};
  end
endmodule
module Memory_198(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_0.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_199(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_1.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_200(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_2.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_201(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_3.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_202(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_4.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_203(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_5.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_204(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_6.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module Memory_205(
  input         clock,
  input  [8:0]  io_address,
  output [31:0] io_dataRead
);
  wire  RamInitSpWf_clk; // @[Memory.scala 65:26]
  wire  RamInitSpWf_we; // @[Memory.scala 65:26]
  wire  RamInitSpWf_en; // @[Memory.scala 65:26]
  wire [8:0] RamInitSpWf_addr; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_di; // @[Memory.scala 65:26]
  wire [31:0] RamInitSpWf_dout; // @[Memory.scala 65:26]
  RamInitSpWf #(.ADDR_WIDTH(9), .DATA_WIDTH(32), .LOAD_FILE("memory_init/tone_init_7.mem")) RamInitSpWf ( // @[Memory.scala 65:26]
    .clk(RamInitSpWf_clk),
    .we(RamInitSpWf_we),
    .en(RamInitSpWf_en),
    .addr(RamInitSpWf_addr),
    .di(RamInitSpWf_di),
    .dout(RamInitSpWf_dout)
  );
  assign io_dataRead = RamInitSpWf_dout; // @[Memory.scala 71:17]
  assign RamInitSpWf_clk = clock; // @[Memory.scala 66:21]
  assign RamInitSpWf_we = 1'h0; // @[Memory.scala 67:20]
  assign RamInitSpWf_en = 1'h1; // @[Memory.scala 68:20]
  assign RamInitSpWf_addr = io_address; // @[Memory.scala 69:22]
  assign RamInitSpWf_di = 32'h0; // @[Memory.scala 70:20]
endmodule
module SoundEngine(
  input        clock,
  input        reset,
  output       io_output_0,
  input  [3:0] io_input
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire  tone_0_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_0_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_0_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_1_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_1_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_1_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_2_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_2_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_2_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_3_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_3_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_3_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_4_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_4_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_4_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_5_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_5_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_5_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_6_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_6_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_6_io_dataRead; // @[SoundEngine.scala 36:23]
  wire  tone_7_clock; // @[SoundEngine.scala 36:23]
  wire [8:0] tone_7_io_address; // @[SoundEngine.scala 36:23]
  wire [31:0] tone_7_io_dataRead; // @[SoundEngine.scala 36:23]
  reg  channel_0; // @[SoundEngine.scala 16:30]
  reg  channel_1; // @[SoundEngine.scala 16:30]
  reg  channel_2; // @[SoundEngine.scala 16:30]
  reg  channel_3; // @[SoundEngine.scala 16:30]
  reg  channel_4; // @[SoundEngine.scala 16:30]
  reg  channel_5; // @[SoundEngine.scala 16:30]
  reg  channel_6; // @[SoundEngine.scala 16:30]
  reg  channel_7; // @[SoundEngine.scala 16:30]
  reg [19:0] cntMilliSecond_0; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_1; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_2; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_3; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_4; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_5; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_6; // @[SoundEngine.scala 17:34]
  reg [19:0] cntMilliSecond_7; // @[SoundEngine.scala 17:34]
  reg [19:0] slowCounter_0; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_1; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_2; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_3; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_4; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_5; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_6; // @[SoundEngine.scala 18:28]
  reg [19:0] slowCounter_7; // @[SoundEngine.scala 18:28]
  reg [31:0] waveCnt_0; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_1; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_2; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_3; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_4; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_5; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_6; // @[SoundEngine.scala 19:28]
  reg [31:0] waveCnt_7; // @[SoundEngine.scala 19:28]
  reg [8:0] toneIndex_0; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_1; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_2; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_3; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_4; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_5; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_6; // @[SoundEngine.scala 20:28]
  reg [8:0] toneIndex_7; // @[SoundEngine.scala 20:28]
  reg  songPlaying_0; // @[SoundEngine.scala 21:28]
  reg  songPlaying_1; // @[SoundEngine.scala 21:28]
  reg  songPlaying_2; // @[SoundEngine.scala 21:28]
  reg  songPlaying_3; // @[SoundEngine.scala 21:28]
  reg  songPlaying_4; // @[SoundEngine.scala 21:28]
  reg  songPlaying_5; // @[SoundEngine.scala 21:28]
  reg  songPlaying_6; // @[SoundEngine.scala 21:28]
  reg  songPlaying_7; // @[SoundEngine.scala 21:28]
  wire  _T_9 = io_input > 4'h0; // @[SoundEngine.scala 27:17]
  wire  _T_10 = io_input <= 4'h8; // @[SoundEngine.scala 27:35]
  wire  _T_11 = _T_9 & _T_10; // @[SoundEngine.scala 27:23]
  wire [3:0] _T_13 = io_input - 4'h1; // @[SoundEngine.scala 28:25]
  wire  _GEN_152 = 3'h0 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_8 = _GEN_152 | songPlaying_0; // @[SoundEngine.scala 28:31]
  wire  _GEN_153 = 3'h1 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_9 = _GEN_153 | songPlaying_1; // @[SoundEngine.scala 28:31]
  wire  _GEN_154 = 3'h2 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_10 = _GEN_154 | songPlaying_2; // @[SoundEngine.scala 28:31]
  wire  _GEN_155 = 3'h3 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_11 = _GEN_155 | songPlaying_3; // @[SoundEngine.scala 28:31]
  wire  _GEN_156 = 3'h4 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_12 = _GEN_156 | songPlaying_4; // @[SoundEngine.scala 28:31]
  wire  _GEN_157 = 3'h5 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_13 = _GEN_157 | songPlaying_5; // @[SoundEngine.scala 28:31]
  wire  _GEN_158 = 3'h6 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_14 = _GEN_158 | songPlaying_6; // @[SoundEngine.scala 28:31]
  wire  _GEN_159 = 3'h7 == _T_13[2:0]; // @[SoundEngine.scala 28:31]
  wire  _GEN_15 = _GEN_159 | songPlaying_7; // @[SoundEngine.scala 28:31]
  reg [19:0] freqReg_0; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_1; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_2; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_3; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_4; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_5; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_6; // @[SoundEngine.scala 49:24]
  reg [19:0] freqReg_7; // @[SoundEngine.scala 49:24]
  reg [11:0] durReg_0; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_1; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_2; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_3; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_4; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_5; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_6; // @[SoundEngine.scala 50:24]
  reg [11:0] durReg_7; // @[SoundEngine.scala 50:24]
  wire  _T_39 = ~songPlaying_0; // @[SoundEngine.scala 56:25]
  wire  _T_40 = slowCounter_0 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_42 = cntMilliSecond_0 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_44 = slowCounter_0 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_45 = freqReg_0 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_47 = waveCnt_0 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_160 = {{12'd0}, freqReg_0}; // @[SoundEngine.scala 81:23]
  wire  _T_48 = waveCnt_0 >= _GEN_160; // @[SoundEngine.scala 81:23]
  wire  _T_49 = ~channel_0; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_161 = {{8'd0}, durReg_0}; // @[SoundEngine.scala 88:28]
  wire  _T_50 = cntMilliSecond_0 >= _GEN_161; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_52 = toneIndex_0 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_53 = durReg_0 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_54 = ~songPlaying_1; // @[SoundEngine.scala 56:25]
  wire  _T_55 = slowCounter_1 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_57 = cntMilliSecond_1 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_59 = slowCounter_1 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_60 = freqReg_1 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_62 = waveCnt_1 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_162 = {{12'd0}, freqReg_1}; // @[SoundEngine.scala 81:23]
  wire  _T_63 = waveCnt_1 >= _GEN_162; // @[SoundEngine.scala 81:23]
  wire  _T_64 = ~channel_1; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_163 = {{8'd0}, durReg_1}; // @[SoundEngine.scala 88:28]
  wire  _T_65 = cntMilliSecond_1 >= _GEN_163; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_67 = toneIndex_1 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_68 = durReg_1 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_69 = ~songPlaying_2; // @[SoundEngine.scala 56:25]
  wire  _T_70 = slowCounter_2 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_72 = cntMilliSecond_2 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_74 = slowCounter_2 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_75 = freqReg_2 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_77 = waveCnt_2 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_164 = {{12'd0}, freqReg_2}; // @[SoundEngine.scala 81:23]
  wire  _T_78 = waveCnt_2 >= _GEN_164; // @[SoundEngine.scala 81:23]
  wire  _T_79 = ~channel_2; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_165 = {{8'd0}, durReg_2}; // @[SoundEngine.scala 88:28]
  wire  _T_80 = cntMilliSecond_2 >= _GEN_165; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_82 = toneIndex_2 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_83 = durReg_2 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_84 = ~songPlaying_3; // @[SoundEngine.scala 56:25]
  wire  _T_85 = slowCounter_3 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_87 = cntMilliSecond_3 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_89 = slowCounter_3 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_90 = freqReg_3 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_92 = waveCnt_3 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_166 = {{12'd0}, freqReg_3}; // @[SoundEngine.scala 81:23]
  wire  _T_93 = waveCnt_3 >= _GEN_166; // @[SoundEngine.scala 81:23]
  wire  _T_94 = ~channel_3; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_167 = {{8'd0}, durReg_3}; // @[SoundEngine.scala 88:28]
  wire  _T_95 = cntMilliSecond_3 >= _GEN_167; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_97 = toneIndex_3 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_98 = durReg_3 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_99 = ~songPlaying_4; // @[SoundEngine.scala 56:25]
  wire  _T_100 = slowCounter_4 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_102 = cntMilliSecond_4 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_104 = slowCounter_4 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_105 = freqReg_4 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_107 = waveCnt_4 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_168 = {{12'd0}, freqReg_4}; // @[SoundEngine.scala 81:23]
  wire  _T_108 = waveCnt_4 >= _GEN_168; // @[SoundEngine.scala 81:23]
  wire  _T_109 = ~channel_4; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_169 = {{8'd0}, durReg_4}; // @[SoundEngine.scala 88:28]
  wire  _T_110 = cntMilliSecond_4 >= _GEN_169; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_112 = toneIndex_4 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_113 = durReg_4 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_114 = ~songPlaying_5; // @[SoundEngine.scala 56:25]
  wire  _T_115 = slowCounter_5 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_117 = cntMilliSecond_5 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_119 = slowCounter_5 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_120 = freqReg_5 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_122 = waveCnt_5 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_170 = {{12'd0}, freqReg_5}; // @[SoundEngine.scala 81:23]
  wire  _T_123 = waveCnt_5 >= _GEN_170; // @[SoundEngine.scala 81:23]
  wire  _T_124 = ~channel_5; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_171 = {{8'd0}, durReg_5}; // @[SoundEngine.scala 88:28]
  wire  _T_125 = cntMilliSecond_5 >= _GEN_171; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_127 = toneIndex_5 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_128 = durReg_5 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_129 = ~songPlaying_6; // @[SoundEngine.scala 56:25]
  wire  _T_130 = slowCounter_6 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_132 = cntMilliSecond_6 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_134 = slowCounter_6 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_135 = freqReg_6 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_137 = waveCnt_6 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_172 = {{12'd0}, freqReg_6}; // @[SoundEngine.scala 81:23]
  wire  _T_138 = waveCnt_6 >= _GEN_172; // @[SoundEngine.scala 81:23]
  wire  _T_139 = ~channel_6; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_173 = {{8'd0}, durReg_6}; // @[SoundEngine.scala 88:28]
  wire  _T_140 = cntMilliSecond_6 >= _GEN_173; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_142 = toneIndex_6 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_143 = durReg_6 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_144 = ~songPlaying_7; // @[SoundEngine.scala 56:25]
  wire  _T_145 = slowCounter_7 == 20'h186a0; // @[SoundEngine.scala 66:25]
  wire [19:0] _T_147 = cntMilliSecond_7 + 20'h1; // @[SoundEngine.scala 68:46]
  wire [19:0] _T_149 = slowCounter_7 + 20'h1; // @[SoundEngine.scala 70:40]
  wire  _T_150 = freqReg_7 == 20'h0; // @[SoundEngine.scala 76:21]
  wire [31:0] _T_152 = waveCnt_7 + 32'h1; // @[SoundEngine.scala 80:32]
  wire [31:0] _GEN_174 = {{12'd0}, freqReg_7}; // @[SoundEngine.scala 81:23]
  wire  _T_153 = waveCnt_7 >= _GEN_174; // @[SoundEngine.scala 81:23]
  wire  _T_154 = ~channel_7; // @[SoundEngine.scala 83:23]
  wire [19:0] _GEN_175 = {{8'd0}, durReg_7}; // @[SoundEngine.scala 88:28]
  wire  _T_155 = cntMilliSecond_7 >= _GEN_175; // @[SoundEngine.scala 88:28]
  wire [8:0] _T_157 = toneIndex_7 + 9'h1; // @[SoundEngine.scala 90:36]
  wire  _T_158 = durReg_7 == 12'hfff; // @[SoundEngine.scala 93:20]
  wire  _T_159 = channel_0 | channel_1; // @[SoundEngine.scala 98:35]
  wire  _T_160 = _T_159 | channel_2; // @[SoundEngine.scala 98:35]
  wire  _T_161 = _T_160 | channel_3; // @[SoundEngine.scala 98:35]
  wire  _T_162 = _T_161 | channel_4; // @[SoundEngine.scala 98:35]
  wire  _T_163 = _T_162 | channel_5; // @[SoundEngine.scala 98:35]
  wire  _T_164 = _T_163 | channel_6; // @[SoundEngine.scala 98:35]
  Memory_198 tone_0 ( // @[SoundEngine.scala 36:23]
    .clock(tone_0_clock),
    .io_address(tone_0_io_address),
    .io_dataRead(tone_0_io_dataRead)
  );
  Memory_199 tone_1 ( // @[SoundEngine.scala 36:23]
    .clock(tone_1_clock),
    .io_address(tone_1_io_address),
    .io_dataRead(tone_1_io_dataRead)
  );
  Memory_200 tone_2 ( // @[SoundEngine.scala 36:23]
    .clock(tone_2_clock),
    .io_address(tone_2_io_address),
    .io_dataRead(tone_2_io_dataRead)
  );
  Memory_201 tone_3 ( // @[SoundEngine.scala 36:23]
    .clock(tone_3_clock),
    .io_address(tone_3_io_address),
    .io_dataRead(tone_3_io_dataRead)
  );
  Memory_202 tone_4 ( // @[SoundEngine.scala 36:23]
    .clock(tone_4_clock),
    .io_address(tone_4_io_address),
    .io_dataRead(tone_4_io_dataRead)
  );
  Memory_203 tone_5 ( // @[SoundEngine.scala 36:23]
    .clock(tone_5_clock),
    .io_address(tone_5_io_address),
    .io_dataRead(tone_5_io_dataRead)
  );
  Memory_204 tone_6 ( // @[SoundEngine.scala 36:23]
    .clock(tone_6_clock),
    .io_address(tone_6_io_address),
    .io_dataRead(tone_6_io_dataRead)
  );
  Memory_205 tone_7 ( // @[SoundEngine.scala 36:23]
    .clock(tone_7_clock),
    .io_address(tone_7_io_address),
    .io_dataRead(tone_7_io_dataRead)
  );
  assign io_output_0 = _T_164 | channel_7; // @[SoundEngine.scala 98:16]
  assign tone_0_clock = clock;
  assign tone_0_io_address = toneIndex_0; // @[SoundEngine.scala 45:24]
  assign tone_1_clock = clock;
  assign tone_1_io_address = toneIndex_1; // @[SoundEngine.scala 45:24]
  assign tone_2_clock = clock;
  assign tone_2_io_address = toneIndex_2; // @[SoundEngine.scala 45:24]
  assign tone_3_clock = clock;
  assign tone_3_io_address = toneIndex_3; // @[SoundEngine.scala 45:24]
  assign tone_4_clock = clock;
  assign tone_4_io_address = toneIndex_4; // @[SoundEngine.scala 45:24]
  assign tone_5_clock = clock;
  assign tone_5_io_address = toneIndex_5; // @[SoundEngine.scala 45:24]
  assign tone_6_clock = clock;
  assign tone_6_io_address = toneIndex_6; // @[SoundEngine.scala 45:24]
  assign tone_7_clock = clock;
  assign tone_7_io_address = toneIndex_7; // @[SoundEngine.scala 45:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  channel_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  channel_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  channel_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  channel_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  channel_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  channel_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  channel_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  channel_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cntMilliSecond_0 = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  cntMilliSecond_1 = _RAND_9[19:0];
  _RAND_10 = {1{`RANDOM}};
  cntMilliSecond_2 = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  cntMilliSecond_3 = _RAND_11[19:0];
  _RAND_12 = {1{`RANDOM}};
  cntMilliSecond_4 = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  cntMilliSecond_5 = _RAND_13[19:0];
  _RAND_14 = {1{`RANDOM}};
  cntMilliSecond_6 = _RAND_14[19:0];
  _RAND_15 = {1{`RANDOM}};
  cntMilliSecond_7 = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  slowCounter_0 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  slowCounter_1 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  slowCounter_2 = _RAND_18[19:0];
  _RAND_19 = {1{`RANDOM}};
  slowCounter_3 = _RAND_19[19:0];
  _RAND_20 = {1{`RANDOM}};
  slowCounter_4 = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  slowCounter_5 = _RAND_21[19:0];
  _RAND_22 = {1{`RANDOM}};
  slowCounter_6 = _RAND_22[19:0];
  _RAND_23 = {1{`RANDOM}};
  slowCounter_7 = _RAND_23[19:0];
  _RAND_24 = {1{`RANDOM}};
  waveCnt_0 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  waveCnt_1 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  waveCnt_2 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  waveCnt_3 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  waveCnt_4 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  waveCnt_5 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  waveCnt_6 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  waveCnt_7 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  toneIndex_0 = _RAND_32[8:0];
  _RAND_33 = {1{`RANDOM}};
  toneIndex_1 = _RAND_33[8:0];
  _RAND_34 = {1{`RANDOM}};
  toneIndex_2 = _RAND_34[8:0];
  _RAND_35 = {1{`RANDOM}};
  toneIndex_3 = _RAND_35[8:0];
  _RAND_36 = {1{`RANDOM}};
  toneIndex_4 = _RAND_36[8:0];
  _RAND_37 = {1{`RANDOM}};
  toneIndex_5 = _RAND_37[8:0];
  _RAND_38 = {1{`RANDOM}};
  toneIndex_6 = _RAND_38[8:0];
  _RAND_39 = {1{`RANDOM}};
  toneIndex_7 = _RAND_39[8:0];
  _RAND_40 = {1{`RANDOM}};
  songPlaying_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  songPlaying_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  songPlaying_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  songPlaying_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  songPlaying_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  songPlaying_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  songPlaying_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  songPlaying_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  freqReg_0 = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  freqReg_1 = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  freqReg_2 = _RAND_50[19:0];
  _RAND_51 = {1{`RANDOM}};
  freqReg_3 = _RAND_51[19:0];
  _RAND_52 = {1{`RANDOM}};
  freqReg_4 = _RAND_52[19:0];
  _RAND_53 = {1{`RANDOM}};
  freqReg_5 = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  freqReg_6 = _RAND_54[19:0];
  _RAND_55 = {1{`RANDOM}};
  freqReg_7 = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  durReg_0 = _RAND_56[11:0];
  _RAND_57 = {1{`RANDOM}};
  durReg_1 = _RAND_57[11:0];
  _RAND_58 = {1{`RANDOM}};
  durReg_2 = _RAND_58[11:0];
  _RAND_59 = {1{`RANDOM}};
  durReg_3 = _RAND_59[11:0];
  _RAND_60 = {1{`RANDOM}};
  durReg_4 = _RAND_60[11:0];
  _RAND_61 = {1{`RANDOM}};
  durReg_5 = _RAND_61[11:0];
  _RAND_62 = {1{`RANDOM}};
  durReg_6 = _RAND_62[11:0];
  _RAND_63 = {1{`RANDOM}};
  durReg_7 = _RAND_63[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      channel_0 <= 1'h0;
    end else if (_T_45) begin
      channel_0 <= 1'h0;
    end else if (_T_48) begin
      channel_0 <= _T_49;
    end else if (_T_39) begin
      channel_0 <= 1'h0;
    end
    if (reset) begin
      channel_1 <= 1'h0;
    end else if (_T_60) begin
      channel_1 <= 1'h0;
    end else if (_T_63) begin
      channel_1 <= _T_64;
    end else if (_T_54) begin
      channel_1 <= 1'h0;
    end
    if (reset) begin
      channel_2 <= 1'h0;
    end else if (_T_75) begin
      channel_2 <= 1'h0;
    end else if (_T_78) begin
      channel_2 <= _T_79;
    end else if (_T_69) begin
      channel_2 <= 1'h0;
    end
    if (reset) begin
      channel_3 <= 1'h0;
    end else if (_T_90) begin
      channel_3 <= 1'h0;
    end else if (_T_93) begin
      channel_3 <= _T_94;
    end else if (_T_84) begin
      channel_3 <= 1'h0;
    end
    if (reset) begin
      channel_4 <= 1'h0;
    end else if (_T_105) begin
      channel_4 <= 1'h0;
    end else if (_T_108) begin
      channel_4 <= _T_109;
    end else if (_T_99) begin
      channel_4 <= 1'h0;
    end
    if (reset) begin
      channel_5 <= 1'h0;
    end else if (_T_120) begin
      channel_5 <= 1'h0;
    end else if (_T_123) begin
      channel_5 <= _T_124;
    end else if (_T_114) begin
      channel_5 <= 1'h0;
    end
    if (reset) begin
      channel_6 <= 1'h0;
    end else if (_T_135) begin
      channel_6 <= 1'h0;
    end else if (_T_138) begin
      channel_6 <= _T_139;
    end else if (_T_129) begin
      channel_6 <= 1'h0;
    end
    if (reset) begin
      channel_7 <= 1'h0;
    end else if (_T_150) begin
      channel_7 <= 1'h0;
    end else if (_T_153) begin
      channel_7 <= _T_154;
    end else if (_T_144) begin
      channel_7 <= 1'h0;
    end
    if (reset) begin
      cntMilliSecond_0 <= 20'h0;
    end else if (_T_50) begin
      cntMilliSecond_0 <= 20'h0;
    end else if (_T_40) begin
      cntMilliSecond_0 <= _T_42;
    end else if (_T_39) begin
      cntMilliSecond_0 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_1 <= 20'h0;
    end else if (_T_65) begin
      cntMilliSecond_1 <= 20'h0;
    end else if (_T_55) begin
      cntMilliSecond_1 <= _T_57;
    end else if (_T_54) begin
      cntMilliSecond_1 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_2 <= 20'h0;
    end else if (_T_80) begin
      cntMilliSecond_2 <= 20'h0;
    end else if (_T_70) begin
      cntMilliSecond_2 <= _T_72;
    end else if (_T_69) begin
      cntMilliSecond_2 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_3 <= 20'h0;
    end else if (_T_95) begin
      cntMilliSecond_3 <= 20'h0;
    end else if (_T_85) begin
      cntMilliSecond_3 <= _T_87;
    end else if (_T_84) begin
      cntMilliSecond_3 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_4 <= 20'h0;
    end else if (_T_110) begin
      cntMilliSecond_4 <= 20'h0;
    end else if (_T_100) begin
      cntMilliSecond_4 <= _T_102;
    end else if (_T_99) begin
      cntMilliSecond_4 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_5 <= 20'h0;
    end else if (_T_125) begin
      cntMilliSecond_5 <= 20'h0;
    end else if (_T_115) begin
      cntMilliSecond_5 <= _T_117;
    end else if (_T_114) begin
      cntMilliSecond_5 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_6 <= 20'h0;
    end else if (_T_140) begin
      cntMilliSecond_6 <= 20'h0;
    end else if (_T_130) begin
      cntMilliSecond_6 <= _T_132;
    end else if (_T_129) begin
      cntMilliSecond_6 <= 20'h0;
    end
    if (reset) begin
      cntMilliSecond_7 <= 20'h0;
    end else if (_T_155) begin
      cntMilliSecond_7 <= 20'h0;
    end else if (_T_145) begin
      cntMilliSecond_7 <= _T_147;
    end else if (_T_144) begin
      cntMilliSecond_7 <= 20'h0;
    end
    if (reset) begin
      slowCounter_0 <= 20'h0;
    end else if (_T_40) begin
      slowCounter_0 <= 20'h0;
    end else begin
      slowCounter_0 <= _T_44;
    end
    if (reset) begin
      slowCounter_1 <= 20'h0;
    end else if (_T_55) begin
      slowCounter_1 <= 20'h0;
    end else begin
      slowCounter_1 <= _T_59;
    end
    if (reset) begin
      slowCounter_2 <= 20'h0;
    end else if (_T_70) begin
      slowCounter_2 <= 20'h0;
    end else begin
      slowCounter_2 <= _T_74;
    end
    if (reset) begin
      slowCounter_3 <= 20'h0;
    end else if (_T_85) begin
      slowCounter_3 <= 20'h0;
    end else begin
      slowCounter_3 <= _T_89;
    end
    if (reset) begin
      slowCounter_4 <= 20'h0;
    end else if (_T_100) begin
      slowCounter_4 <= 20'h0;
    end else begin
      slowCounter_4 <= _T_104;
    end
    if (reset) begin
      slowCounter_5 <= 20'h0;
    end else if (_T_115) begin
      slowCounter_5 <= 20'h0;
    end else begin
      slowCounter_5 <= _T_119;
    end
    if (reset) begin
      slowCounter_6 <= 20'h0;
    end else if (_T_130) begin
      slowCounter_6 <= 20'h0;
    end else begin
      slowCounter_6 <= _T_134;
    end
    if (reset) begin
      slowCounter_7 <= 20'h0;
    end else if (_T_145) begin
      slowCounter_7 <= 20'h0;
    end else begin
      slowCounter_7 <= _T_149;
    end
    if (reset) begin
      waveCnt_0 <= 32'h0;
    end else if (_T_45) begin
      waveCnt_0 <= 32'h0;
    end else if (_T_48) begin
      waveCnt_0 <= 32'h0;
    end else begin
      waveCnt_0 <= _T_47;
    end
    if (reset) begin
      waveCnt_1 <= 32'h0;
    end else if (_T_60) begin
      waveCnt_1 <= 32'h0;
    end else if (_T_63) begin
      waveCnt_1 <= 32'h0;
    end else begin
      waveCnt_1 <= _T_62;
    end
    if (reset) begin
      waveCnt_2 <= 32'h0;
    end else if (_T_75) begin
      waveCnt_2 <= 32'h0;
    end else if (_T_78) begin
      waveCnt_2 <= 32'h0;
    end else begin
      waveCnt_2 <= _T_77;
    end
    if (reset) begin
      waveCnt_3 <= 32'h0;
    end else if (_T_90) begin
      waveCnt_3 <= 32'h0;
    end else if (_T_93) begin
      waveCnt_3 <= 32'h0;
    end else begin
      waveCnt_3 <= _T_92;
    end
    if (reset) begin
      waveCnt_4 <= 32'h0;
    end else if (_T_105) begin
      waveCnt_4 <= 32'h0;
    end else if (_T_108) begin
      waveCnt_4 <= 32'h0;
    end else begin
      waveCnt_4 <= _T_107;
    end
    if (reset) begin
      waveCnt_5 <= 32'h0;
    end else if (_T_120) begin
      waveCnt_5 <= 32'h0;
    end else if (_T_123) begin
      waveCnt_5 <= 32'h0;
    end else begin
      waveCnt_5 <= _T_122;
    end
    if (reset) begin
      waveCnt_6 <= 32'h0;
    end else if (_T_135) begin
      waveCnt_6 <= 32'h0;
    end else if (_T_138) begin
      waveCnt_6 <= 32'h0;
    end else begin
      waveCnt_6 <= _T_137;
    end
    if (reset) begin
      waveCnt_7 <= 32'h0;
    end else if (_T_150) begin
      waveCnt_7 <= 32'h0;
    end else if (_T_153) begin
      waveCnt_7 <= 32'h0;
    end else begin
      waveCnt_7 <= _T_152;
    end
    if (reset) begin
      toneIndex_0 <= 9'h0;
    end else if (_T_50) begin
      toneIndex_0 <= _T_52;
    end else if (_T_39) begin
      toneIndex_0 <= 9'h0;
    end
    if (reset) begin
      toneIndex_1 <= 9'h0;
    end else if (_T_65) begin
      toneIndex_1 <= _T_67;
    end else if (_T_54) begin
      toneIndex_1 <= 9'h0;
    end
    if (reset) begin
      toneIndex_2 <= 9'h0;
    end else if (_T_80) begin
      toneIndex_2 <= _T_82;
    end else if (_T_69) begin
      toneIndex_2 <= 9'h0;
    end
    if (reset) begin
      toneIndex_3 <= 9'h0;
    end else if (_T_95) begin
      toneIndex_3 <= _T_97;
    end else if (_T_84) begin
      toneIndex_3 <= 9'h0;
    end
    if (reset) begin
      toneIndex_4 <= 9'h0;
    end else if (_T_110) begin
      toneIndex_4 <= _T_112;
    end else if (_T_99) begin
      toneIndex_4 <= 9'h0;
    end
    if (reset) begin
      toneIndex_5 <= 9'h0;
    end else if (_T_125) begin
      toneIndex_5 <= _T_127;
    end else if (_T_114) begin
      toneIndex_5 <= 9'h0;
    end
    if (reset) begin
      toneIndex_6 <= 9'h0;
    end else if (_T_140) begin
      toneIndex_6 <= _T_142;
    end else if (_T_129) begin
      toneIndex_6 <= 9'h0;
    end
    if (reset) begin
      toneIndex_7 <= 9'h0;
    end else if (_T_155) begin
      toneIndex_7 <= _T_157;
    end else if (_T_144) begin
      toneIndex_7 <= 9'h0;
    end
    if (reset) begin
      songPlaying_0 <= 1'h0;
    end else if (_T_53) begin
      songPlaying_0 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_0 <= _GEN_8;
    end
    if (reset) begin
      songPlaying_1 <= 1'h0;
    end else if (_T_68) begin
      songPlaying_1 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_1 <= _GEN_9;
    end
    if (reset) begin
      songPlaying_2 <= 1'h0;
    end else if (_T_83) begin
      songPlaying_2 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_2 <= _GEN_10;
    end
    if (reset) begin
      songPlaying_3 <= 1'h0;
    end else if (_T_98) begin
      songPlaying_3 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_3 <= _GEN_11;
    end
    if (reset) begin
      songPlaying_4 <= 1'h0;
    end else if (_T_113) begin
      songPlaying_4 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_4 <= _GEN_12;
    end
    if (reset) begin
      songPlaying_5 <= 1'h0;
    end else if (_T_128) begin
      songPlaying_5 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_5 <= _GEN_13;
    end
    if (reset) begin
      songPlaying_6 <= 1'h0;
    end else if (_T_143) begin
      songPlaying_6 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_6 <= _GEN_14;
    end
    if (reset) begin
      songPlaying_7 <= 1'h0;
    end else if (_T_158) begin
      songPlaying_7 <= 1'h0;
    end else if (_T_11) begin
      songPlaying_7 <= _GEN_15;
    end
    freqReg_0 <= tone_0_io_dataRead[31:12];
    freqReg_1 <= tone_1_io_dataRead[31:12];
    freqReg_2 <= tone_2_io_dataRead[31:12];
    freqReg_3 <= tone_3_io_dataRead[31:12];
    freqReg_4 <= tone_4_io_dataRead[31:12];
    freqReg_5 <= tone_5_io_dataRead[31:12];
    freqReg_6 <= tone_6_io_dataRead[31:12];
    freqReg_7 <= tone_7_io_dataRead[31:12];
    durReg_0 <= tone_0_io_dataRead[11:0];
    durReg_1 <= tone_1_io_dataRead[11:0];
    durReg_2 <= tone_2_io_dataRead[11:0];
    durReg_3 <= tone_3_io_dataRead[11:0];
    durReg_4 <= tone_4_io_dataRead[11:0];
    durReg_5 <= tone_5_io_dataRead[11:0];
    durReg_6 <= tone_6_io_dataRead[11:0];
    durReg_7 <= tone_7_io_dataRead[11:0];
  end
endmodule
module BoxDetection(
  input         clock,
  input  [10:0] io_boxXPosition_0,
  input  [10:0] io_boxXPosition_2,
  input  [10:0] io_boxXPosition_3,
  input  [10:0] io_boxXPosition_4,
  input  [10:0] io_boxXPosition_5,
  input  [10:0] io_boxXPosition_6,
  input  [10:0] io_boxXPosition_7,
  input  [10:0] io_boxXPosition_8,
  input  [10:0] io_boxXPosition_9,
  input  [10:0] io_boxXPosition_10,
  input  [10:0] io_boxXPosition_11,
  input  [10:0] io_boxXPosition_12,
  input  [10:0] io_boxXPosition_13,
  input  [10:0] io_boxXPosition_14,
  input  [10:0] io_boxXPosition_15,
  input  [10:0] io_boxXPosition_16,
  input  [10:0] io_boxXPosition_17,
  input  [9:0]  io_boxYPosition_0,
  input  [9:0]  io_boxYPosition_2,
  input  [9:0]  io_boxYPosition_3,
  input  [9:0]  io_boxYPosition_4,
  input  [9:0]  io_boxYPosition_5,
  input  [9:0]  io_boxYPosition_6,
  input  [9:0]  io_boxYPosition_7,
  input  [9:0]  io_boxYPosition_8,
  input  [9:0]  io_boxYPosition_9,
  input  [9:0]  io_boxYPosition_10,
  input  [9:0]  io_boxYPosition_11,
  input  [9:0]  io_boxYPosition_12,
  input  [9:0]  io_boxYPosition_13,
  input  [9:0]  io_boxYPosition_14,
  input  [9:0]  io_boxYPosition_15,
  input  [9:0]  io_boxYPosition_16,
  input  [9:0]  io_boxYPosition_17,
  output        io_overlap_0_7,
  output        io_overlap_0_8,
  output        io_overlap_0_9,
  output        io_overlap_0_10,
  output        io_overlap_0_11,
  output        io_overlap_0_12,
  output        io_overlap_0_13,
  output        io_overlap_0_14,
  output        io_overlap_0_15,
  output        io_overlap_0_16,
  output        io_overlap_0_17,
  output        io_overlap_2_7,
  output        io_overlap_2_8,
  output        io_overlap_2_9,
  output        io_overlap_2_10,
  output        io_overlap_2_11,
  output        io_overlap_2_12,
  output        io_overlap_2_13,
  output        io_overlap_2_14,
  output        io_overlap_2_15,
  output        io_overlap_2_16,
  output        io_overlap_2_17,
  output        io_overlap_3_7,
  output        io_overlap_3_8,
  output        io_overlap_3_9,
  output        io_overlap_3_10,
  output        io_overlap_3_11,
  output        io_overlap_3_12,
  output        io_overlap_3_13,
  output        io_overlap_3_14,
  output        io_overlap_3_15,
  output        io_overlap_3_16,
  output        io_overlap_3_17,
  output        io_overlap_4_7,
  output        io_overlap_4_8,
  output        io_overlap_4_9,
  output        io_overlap_4_10,
  output        io_overlap_4_11,
  output        io_overlap_4_12,
  output        io_overlap_4_13,
  output        io_overlap_4_14,
  output        io_overlap_4_15,
  output        io_overlap_4_16,
  output        io_overlap_4_17,
  output        io_overlap_5_7,
  output        io_overlap_5_8,
  output        io_overlap_5_9,
  output        io_overlap_5_10,
  output        io_overlap_5_11,
  output        io_overlap_5_12,
  output        io_overlap_5_13,
  output        io_overlap_5_14,
  output        io_overlap_5_15,
  output        io_overlap_5_16,
  output        io_overlap_5_17,
  output        io_overlap_6_7,
  output        io_overlap_6_8,
  output        io_overlap_6_9,
  output        io_overlap_6_10,
  output        io_overlap_6_11,
  output        io_overlap_6_12,
  output        io_overlap_6_13,
  output        io_overlap_6_14,
  output        io_overlap_6_15,
  output        io_overlap_6_17
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
`endif // RANDOMIZE_REG_INIT
  wire [10:0] _T_2 = $signed(io_boxXPosition_0) + 11'sh20; // @[BoxDetection.scala 18:36]
  wire [9:0] _T_5 = $signed(io_boxYPosition_0) + 10'sh20; // @[BoxDetection.scala 19:36]
  wire [10:0] _T_34 = $signed(io_boxXPosition_2) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_37 = $signed(io_boxYPosition_2) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_47 = $signed(io_boxXPosition_3) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_50 = $signed(io_boxYPosition_3) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_60 = $signed(io_boxXPosition_4) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_63 = $signed(io_boxYPosition_4) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_73 = $signed(io_boxXPosition_5) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_76 = $signed(io_boxYPosition_5) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_86 = $signed(io_boxXPosition_6) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_89 = $signed(io_boxYPosition_6) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire [10:0] _T_99 = $signed(io_boxXPosition_7) + 11'sh8; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_102 = $signed(io_boxYPosition_7) + 10'sh8; // @[BoxDetection.scala 25:38]
  wire  _T_103 = $signed(io_boxXPosition_0) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_104 = $signed(io_boxXPosition_7) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_105 = _T_103 & _T_104; // @[BoxDetection.scala 27:41]
  wire  _T_106 = $signed(io_boxYPosition_0) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_107 = _T_105 & _T_106; // @[BoxDetection.scala 27:60]
  wire  _T_108 = $signed(io_boxYPosition_7) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_112 = $signed(io_boxXPosition_8) + 11'sh10; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_115 = $signed(io_boxYPosition_8) + 10'sh10; // @[BoxDetection.scala 25:38]
  wire  _T_116 = $signed(io_boxXPosition_0) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_117 = $signed(io_boxXPosition_8) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_118 = _T_116 & _T_117; // @[BoxDetection.scala 27:41]
  wire  _T_119 = $signed(io_boxYPosition_0) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_120 = _T_118 & _T_119; // @[BoxDetection.scala 27:60]
  wire  _T_121 = $signed(io_boxYPosition_8) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_125 = $signed(io_boxXPosition_9) + 11'sh1c; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_128 = $signed(io_boxYPosition_9) + 10'sh1c; // @[BoxDetection.scala 25:38]
  wire  _T_129 = $signed(io_boxXPosition_0) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_130 = $signed(io_boxXPosition_9) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_131 = _T_129 & _T_130; // @[BoxDetection.scala 27:41]
  wire  _T_132 = $signed(io_boxYPosition_0) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_133 = _T_131 & _T_132; // @[BoxDetection.scala 27:60]
  wire  _T_134 = $signed(io_boxYPosition_9) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_138 = $signed(io_boxXPosition_10) + 11'sh1c; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_141 = $signed(io_boxYPosition_10) + 10'sh1c; // @[BoxDetection.scala 25:38]
  wire  _T_142 = $signed(io_boxXPosition_0) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_143 = $signed(io_boxXPosition_10) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_144 = _T_142 & _T_143; // @[BoxDetection.scala 27:41]
  wire  _T_145 = $signed(io_boxYPosition_0) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_146 = _T_144 & _T_145; // @[BoxDetection.scala 27:60]
  wire  _T_147 = $signed(io_boxYPosition_10) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_151 = $signed(io_boxXPosition_11) + 11'sh1c; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_154 = $signed(io_boxYPosition_11) + 10'sh1c; // @[BoxDetection.scala 25:38]
  wire  _T_155 = $signed(io_boxXPosition_0) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_156 = $signed(io_boxXPosition_11) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_157 = _T_155 & _T_156; // @[BoxDetection.scala 27:41]
  wire  _T_158 = $signed(io_boxYPosition_0) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_159 = _T_157 & _T_158; // @[BoxDetection.scala 27:60]
  wire  _T_160 = $signed(io_boxYPosition_11) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_164 = $signed(io_boxXPosition_12) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_167 = $signed(io_boxYPosition_12) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_168 = $signed(io_boxXPosition_0) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_169 = $signed(io_boxXPosition_12) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_170 = _T_168 & _T_169; // @[BoxDetection.scala 27:41]
  wire  _T_171 = $signed(io_boxYPosition_0) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_172 = _T_170 & _T_171; // @[BoxDetection.scala 27:60]
  wire  _T_173 = $signed(io_boxYPosition_12) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_177 = $signed(io_boxXPosition_13) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_180 = $signed(io_boxYPosition_13) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_181 = $signed(io_boxXPosition_0) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_182 = $signed(io_boxXPosition_13) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_183 = _T_181 & _T_182; // @[BoxDetection.scala 27:41]
  wire  _T_184 = $signed(io_boxYPosition_0) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_185 = _T_183 & _T_184; // @[BoxDetection.scala 27:60]
  wire  _T_186 = $signed(io_boxYPosition_13) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_190 = $signed(io_boxXPosition_14) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_193 = $signed(io_boxYPosition_14) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_194 = $signed(io_boxXPosition_0) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_195 = $signed(io_boxXPosition_14) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_196 = _T_194 & _T_195; // @[BoxDetection.scala 27:41]
  wire  _T_197 = $signed(io_boxYPosition_0) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_198 = _T_196 & _T_197; // @[BoxDetection.scala 27:60]
  wire  _T_199 = $signed(io_boxYPosition_14) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_203 = $signed(io_boxXPosition_15) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_206 = $signed(io_boxYPosition_15) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_207 = $signed(io_boxXPosition_0) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_208 = $signed(io_boxXPosition_15) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_209 = _T_207 & _T_208; // @[BoxDetection.scala 27:41]
  wire  _T_210 = $signed(io_boxYPosition_0) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_211 = _T_209 & _T_210; // @[BoxDetection.scala 27:60]
  wire  _T_212 = $signed(io_boxYPosition_15) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_216 = $signed(io_boxXPosition_16) + 11'sh20; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_219 = $signed(io_boxYPosition_16) + 10'sh20; // @[BoxDetection.scala 25:38]
  wire  _T_220 = $signed(io_boxXPosition_0) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_221 = $signed(io_boxXPosition_16) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_222 = _T_220 & _T_221; // @[BoxDetection.scala 27:41]
  wire  _T_223 = $signed(io_boxYPosition_0) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_224 = _T_222 & _T_223; // @[BoxDetection.scala 27:60]
  wire  _T_225 = $signed(io_boxYPosition_16) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire [10:0] _T_229 = $signed(io_boxXPosition_17) + 11'sh60; // @[BoxDetection.scala 24:38]
  wire [9:0] _T_232 = $signed(io_boxYPosition_17) + 10'sh60; // @[BoxDetection.scala 25:38]
  wire  _T_233 = $signed(io_boxXPosition_0) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_234 = $signed(io_boxXPosition_17) < $signed(_T_2); // @[BoxDetection.scala 27:51]
  wire  _T_235 = _T_233 & _T_234; // @[BoxDetection.scala 27:41]
  wire  _T_236 = $signed(io_boxYPosition_0) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_237 = _T_235 & _T_236; // @[BoxDetection.scala 27:60]
  wire  _T_238 = $signed(io_boxYPosition_17) < $signed(_T_5); // @[BoxDetection.scala 28:35]
  wire  _T_583 = $signed(io_boxXPosition_2) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_584 = $signed(io_boxXPosition_7) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_585 = _T_583 & _T_584; // @[BoxDetection.scala 27:41]
  wire  _T_586 = $signed(io_boxYPosition_2) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_587 = _T_585 & _T_586; // @[BoxDetection.scala 27:60]
  wire  _T_588 = $signed(io_boxYPosition_7) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_596 = $signed(io_boxXPosition_2) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_597 = $signed(io_boxXPosition_8) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_598 = _T_596 & _T_597; // @[BoxDetection.scala 27:41]
  wire  _T_599 = $signed(io_boxYPosition_2) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_600 = _T_598 & _T_599; // @[BoxDetection.scala 27:60]
  wire  _T_601 = $signed(io_boxYPosition_8) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_609 = $signed(io_boxXPosition_2) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_610 = $signed(io_boxXPosition_9) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_611 = _T_609 & _T_610; // @[BoxDetection.scala 27:41]
  wire  _T_612 = $signed(io_boxYPosition_2) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_613 = _T_611 & _T_612; // @[BoxDetection.scala 27:60]
  wire  _T_614 = $signed(io_boxYPosition_9) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_622 = $signed(io_boxXPosition_2) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_623 = $signed(io_boxXPosition_10) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_624 = _T_622 & _T_623; // @[BoxDetection.scala 27:41]
  wire  _T_625 = $signed(io_boxYPosition_2) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_626 = _T_624 & _T_625; // @[BoxDetection.scala 27:60]
  wire  _T_627 = $signed(io_boxYPosition_10) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_635 = $signed(io_boxXPosition_2) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_636 = $signed(io_boxXPosition_11) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_637 = _T_635 & _T_636; // @[BoxDetection.scala 27:41]
  wire  _T_638 = $signed(io_boxYPosition_2) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_639 = _T_637 & _T_638; // @[BoxDetection.scala 27:60]
  wire  _T_640 = $signed(io_boxYPosition_11) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_648 = $signed(io_boxXPosition_2) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_649 = $signed(io_boxXPosition_12) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_650 = _T_648 & _T_649; // @[BoxDetection.scala 27:41]
  wire  _T_651 = $signed(io_boxYPosition_2) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_652 = _T_650 & _T_651; // @[BoxDetection.scala 27:60]
  wire  _T_653 = $signed(io_boxYPosition_12) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_661 = $signed(io_boxXPosition_2) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_662 = $signed(io_boxXPosition_13) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_663 = _T_661 & _T_662; // @[BoxDetection.scala 27:41]
  wire  _T_664 = $signed(io_boxYPosition_2) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_665 = _T_663 & _T_664; // @[BoxDetection.scala 27:60]
  wire  _T_666 = $signed(io_boxYPosition_13) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_674 = $signed(io_boxXPosition_2) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_675 = $signed(io_boxXPosition_14) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_676 = _T_674 & _T_675; // @[BoxDetection.scala 27:41]
  wire  _T_677 = $signed(io_boxYPosition_2) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_678 = _T_676 & _T_677; // @[BoxDetection.scala 27:60]
  wire  _T_679 = $signed(io_boxYPosition_14) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_687 = $signed(io_boxXPosition_2) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_688 = $signed(io_boxXPosition_15) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_689 = _T_687 & _T_688; // @[BoxDetection.scala 27:41]
  wire  _T_690 = $signed(io_boxYPosition_2) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_691 = _T_689 & _T_690; // @[BoxDetection.scala 27:60]
  wire  _T_692 = $signed(io_boxYPosition_15) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_700 = $signed(io_boxXPosition_2) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_701 = $signed(io_boxXPosition_16) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_702 = _T_700 & _T_701; // @[BoxDetection.scala 27:41]
  wire  _T_703 = $signed(io_boxYPosition_2) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_704 = _T_702 & _T_703; // @[BoxDetection.scala 27:60]
  wire  _T_705 = $signed(io_boxYPosition_16) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_713 = $signed(io_boxXPosition_2) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_714 = $signed(io_boxXPosition_17) < $signed(_T_34); // @[BoxDetection.scala 27:51]
  wire  _T_715 = _T_713 & _T_714; // @[BoxDetection.scala 27:41]
  wire  _T_716 = $signed(io_boxYPosition_2) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_717 = _T_715 & _T_716; // @[BoxDetection.scala 27:60]
  wire  _T_718 = $signed(io_boxYPosition_17) < $signed(_T_37); // @[BoxDetection.scala 28:35]
  wire  _T_823 = $signed(io_boxXPosition_3) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_824 = $signed(io_boxXPosition_7) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_825 = _T_823 & _T_824; // @[BoxDetection.scala 27:41]
  wire  _T_826 = $signed(io_boxYPosition_3) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_827 = _T_825 & _T_826; // @[BoxDetection.scala 27:60]
  wire  _T_828 = $signed(io_boxYPosition_7) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_836 = $signed(io_boxXPosition_3) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_837 = $signed(io_boxXPosition_8) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_838 = _T_836 & _T_837; // @[BoxDetection.scala 27:41]
  wire  _T_839 = $signed(io_boxYPosition_3) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_840 = _T_838 & _T_839; // @[BoxDetection.scala 27:60]
  wire  _T_841 = $signed(io_boxYPosition_8) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_849 = $signed(io_boxXPosition_3) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_850 = $signed(io_boxXPosition_9) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_851 = _T_849 & _T_850; // @[BoxDetection.scala 27:41]
  wire  _T_852 = $signed(io_boxYPosition_3) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_853 = _T_851 & _T_852; // @[BoxDetection.scala 27:60]
  wire  _T_854 = $signed(io_boxYPosition_9) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_862 = $signed(io_boxXPosition_3) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_863 = $signed(io_boxXPosition_10) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_864 = _T_862 & _T_863; // @[BoxDetection.scala 27:41]
  wire  _T_865 = $signed(io_boxYPosition_3) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_866 = _T_864 & _T_865; // @[BoxDetection.scala 27:60]
  wire  _T_867 = $signed(io_boxYPosition_10) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_875 = $signed(io_boxXPosition_3) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_876 = $signed(io_boxXPosition_11) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_877 = _T_875 & _T_876; // @[BoxDetection.scala 27:41]
  wire  _T_878 = $signed(io_boxYPosition_3) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_879 = _T_877 & _T_878; // @[BoxDetection.scala 27:60]
  wire  _T_880 = $signed(io_boxYPosition_11) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_888 = $signed(io_boxXPosition_3) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_889 = $signed(io_boxXPosition_12) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_890 = _T_888 & _T_889; // @[BoxDetection.scala 27:41]
  wire  _T_891 = $signed(io_boxYPosition_3) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_892 = _T_890 & _T_891; // @[BoxDetection.scala 27:60]
  wire  _T_893 = $signed(io_boxYPosition_12) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_901 = $signed(io_boxXPosition_3) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_902 = $signed(io_boxXPosition_13) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_903 = _T_901 & _T_902; // @[BoxDetection.scala 27:41]
  wire  _T_904 = $signed(io_boxYPosition_3) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_905 = _T_903 & _T_904; // @[BoxDetection.scala 27:60]
  wire  _T_906 = $signed(io_boxYPosition_13) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_914 = $signed(io_boxXPosition_3) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_915 = $signed(io_boxXPosition_14) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_916 = _T_914 & _T_915; // @[BoxDetection.scala 27:41]
  wire  _T_917 = $signed(io_boxYPosition_3) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_918 = _T_916 & _T_917; // @[BoxDetection.scala 27:60]
  wire  _T_919 = $signed(io_boxYPosition_14) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_927 = $signed(io_boxXPosition_3) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_928 = $signed(io_boxXPosition_15) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_929 = _T_927 & _T_928; // @[BoxDetection.scala 27:41]
  wire  _T_930 = $signed(io_boxYPosition_3) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_931 = _T_929 & _T_930; // @[BoxDetection.scala 27:60]
  wire  _T_932 = $signed(io_boxYPosition_15) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_940 = $signed(io_boxXPosition_3) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_941 = $signed(io_boxXPosition_16) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_942 = _T_940 & _T_941; // @[BoxDetection.scala 27:41]
  wire  _T_943 = $signed(io_boxYPosition_3) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_944 = _T_942 & _T_943; // @[BoxDetection.scala 27:60]
  wire  _T_945 = $signed(io_boxYPosition_16) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_953 = $signed(io_boxXPosition_3) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_954 = $signed(io_boxXPosition_17) < $signed(_T_47); // @[BoxDetection.scala 27:51]
  wire  _T_955 = _T_953 & _T_954; // @[BoxDetection.scala 27:41]
  wire  _T_956 = $signed(io_boxYPosition_3) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_957 = _T_955 & _T_956; // @[BoxDetection.scala 27:60]
  wire  _T_958 = $signed(io_boxYPosition_17) < $signed(_T_50); // @[BoxDetection.scala 28:35]
  wire  _T_1063 = $signed(io_boxXPosition_4) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_1064 = $signed(io_boxXPosition_7) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1065 = _T_1063 & _T_1064; // @[BoxDetection.scala 27:41]
  wire  _T_1066 = $signed(io_boxYPosition_4) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_1067 = _T_1065 & _T_1066; // @[BoxDetection.scala 27:60]
  wire  _T_1068 = $signed(io_boxYPosition_7) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1076 = $signed(io_boxXPosition_4) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_1077 = $signed(io_boxXPosition_8) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1078 = _T_1076 & _T_1077; // @[BoxDetection.scala 27:41]
  wire  _T_1079 = $signed(io_boxYPosition_4) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_1080 = _T_1078 & _T_1079; // @[BoxDetection.scala 27:60]
  wire  _T_1081 = $signed(io_boxYPosition_8) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1089 = $signed(io_boxXPosition_4) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_1090 = $signed(io_boxXPosition_9) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1091 = _T_1089 & _T_1090; // @[BoxDetection.scala 27:41]
  wire  _T_1092 = $signed(io_boxYPosition_4) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_1093 = _T_1091 & _T_1092; // @[BoxDetection.scala 27:60]
  wire  _T_1094 = $signed(io_boxYPosition_9) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1102 = $signed(io_boxXPosition_4) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_1103 = $signed(io_boxXPosition_10) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1104 = _T_1102 & _T_1103; // @[BoxDetection.scala 27:41]
  wire  _T_1105 = $signed(io_boxYPosition_4) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_1106 = _T_1104 & _T_1105; // @[BoxDetection.scala 27:60]
  wire  _T_1107 = $signed(io_boxYPosition_10) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1115 = $signed(io_boxXPosition_4) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_1116 = $signed(io_boxXPosition_11) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1117 = _T_1115 & _T_1116; // @[BoxDetection.scala 27:41]
  wire  _T_1118 = $signed(io_boxYPosition_4) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_1119 = _T_1117 & _T_1118; // @[BoxDetection.scala 27:60]
  wire  _T_1120 = $signed(io_boxYPosition_11) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1128 = $signed(io_boxXPosition_4) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_1129 = $signed(io_boxXPosition_12) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1130 = _T_1128 & _T_1129; // @[BoxDetection.scala 27:41]
  wire  _T_1131 = $signed(io_boxYPosition_4) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_1132 = _T_1130 & _T_1131; // @[BoxDetection.scala 27:60]
  wire  _T_1133 = $signed(io_boxYPosition_12) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1141 = $signed(io_boxXPosition_4) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_1142 = $signed(io_boxXPosition_13) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1143 = _T_1141 & _T_1142; // @[BoxDetection.scala 27:41]
  wire  _T_1144 = $signed(io_boxYPosition_4) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_1145 = _T_1143 & _T_1144; // @[BoxDetection.scala 27:60]
  wire  _T_1146 = $signed(io_boxYPosition_13) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1154 = $signed(io_boxXPosition_4) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_1155 = $signed(io_boxXPosition_14) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1156 = _T_1154 & _T_1155; // @[BoxDetection.scala 27:41]
  wire  _T_1157 = $signed(io_boxYPosition_4) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_1158 = _T_1156 & _T_1157; // @[BoxDetection.scala 27:60]
  wire  _T_1159 = $signed(io_boxYPosition_14) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1167 = $signed(io_boxXPosition_4) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_1168 = $signed(io_boxXPosition_15) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1169 = _T_1167 & _T_1168; // @[BoxDetection.scala 27:41]
  wire  _T_1170 = $signed(io_boxYPosition_4) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_1171 = _T_1169 & _T_1170; // @[BoxDetection.scala 27:60]
  wire  _T_1172 = $signed(io_boxYPosition_15) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1180 = $signed(io_boxXPosition_4) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_1181 = $signed(io_boxXPosition_16) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1182 = _T_1180 & _T_1181; // @[BoxDetection.scala 27:41]
  wire  _T_1183 = $signed(io_boxYPosition_4) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_1184 = _T_1182 & _T_1183; // @[BoxDetection.scala 27:60]
  wire  _T_1185 = $signed(io_boxYPosition_16) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1193 = $signed(io_boxXPosition_4) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_1194 = $signed(io_boxXPosition_17) < $signed(_T_60); // @[BoxDetection.scala 27:51]
  wire  _T_1195 = _T_1193 & _T_1194; // @[BoxDetection.scala 27:41]
  wire  _T_1196 = $signed(io_boxYPosition_4) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_1197 = _T_1195 & _T_1196; // @[BoxDetection.scala 27:60]
  wire  _T_1198 = $signed(io_boxYPosition_17) < $signed(_T_63); // @[BoxDetection.scala 28:35]
  wire  _T_1303 = $signed(io_boxXPosition_5) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_1304 = $signed(io_boxXPosition_7) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1305 = _T_1303 & _T_1304; // @[BoxDetection.scala 27:41]
  wire  _T_1306 = $signed(io_boxYPosition_5) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_1307 = _T_1305 & _T_1306; // @[BoxDetection.scala 27:60]
  wire  _T_1308 = $signed(io_boxYPosition_7) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1316 = $signed(io_boxXPosition_5) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_1317 = $signed(io_boxXPosition_8) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1318 = _T_1316 & _T_1317; // @[BoxDetection.scala 27:41]
  wire  _T_1319 = $signed(io_boxYPosition_5) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_1320 = _T_1318 & _T_1319; // @[BoxDetection.scala 27:60]
  wire  _T_1321 = $signed(io_boxYPosition_8) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1329 = $signed(io_boxXPosition_5) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_1330 = $signed(io_boxXPosition_9) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1331 = _T_1329 & _T_1330; // @[BoxDetection.scala 27:41]
  wire  _T_1332 = $signed(io_boxYPosition_5) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_1333 = _T_1331 & _T_1332; // @[BoxDetection.scala 27:60]
  wire  _T_1334 = $signed(io_boxYPosition_9) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1342 = $signed(io_boxXPosition_5) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_1343 = $signed(io_boxXPosition_10) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1344 = _T_1342 & _T_1343; // @[BoxDetection.scala 27:41]
  wire  _T_1345 = $signed(io_boxYPosition_5) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_1346 = _T_1344 & _T_1345; // @[BoxDetection.scala 27:60]
  wire  _T_1347 = $signed(io_boxYPosition_10) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1355 = $signed(io_boxXPosition_5) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_1356 = $signed(io_boxXPosition_11) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1357 = _T_1355 & _T_1356; // @[BoxDetection.scala 27:41]
  wire  _T_1358 = $signed(io_boxYPosition_5) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_1359 = _T_1357 & _T_1358; // @[BoxDetection.scala 27:60]
  wire  _T_1360 = $signed(io_boxYPosition_11) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1368 = $signed(io_boxXPosition_5) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_1369 = $signed(io_boxXPosition_12) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1370 = _T_1368 & _T_1369; // @[BoxDetection.scala 27:41]
  wire  _T_1371 = $signed(io_boxYPosition_5) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_1372 = _T_1370 & _T_1371; // @[BoxDetection.scala 27:60]
  wire  _T_1373 = $signed(io_boxYPosition_12) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1381 = $signed(io_boxXPosition_5) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_1382 = $signed(io_boxXPosition_13) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1383 = _T_1381 & _T_1382; // @[BoxDetection.scala 27:41]
  wire  _T_1384 = $signed(io_boxYPosition_5) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_1385 = _T_1383 & _T_1384; // @[BoxDetection.scala 27:60]
  wire  _T_1386 = $signed(io_boxYPosition_13) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1394 = $signed(io_boxXPosition_5) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_1395 = $signed(io_boxXPosition_14) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1396 = _T_1394 & _T_1395; // @[BoxDetection.scala 27:41]
  wire  _T_1397 = $signed(io_boxYPosition_5) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_1398 = _T_1396 & _T_1397; // @[BoxDetection.scala 27:60]
  wire  _T_1399 = $signed(io_boxYPosition_14) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1407 = $signed(io_boxXPosition_5) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_1408 = $signed(io_boxXPosition_15) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1409 = _T_1407 & _T_1408; // @[BoxDetection.scala 27:41]
  wire  _T_1410 = $signed(io_boxYPosition_5) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_1411 = _T_1409 & _T_1410; // @[BoxDetection.scala 27:60]
  wire  _T_1412 = $signed(io_boxYPosition_15) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1420 = $signed(io_boxXPosition_5) < $signed(_T_216); // @[BoxDetection.scala 27:32]
  wire  _T_1421 = $signed(io_boxXPosition_16) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1422 = _T_1420 & _T_1421; // @[BoxDetection.scala 27:41]
  wire  _T_1423 = $signed(io_boxYPosition_5) < $signed(_T_219); // @[BoxDetection.scala 28:16]
  wire  _T_1424 = _T_1422 & _T_1423; // @[BoxDetection.scala 27:60]
  wire  _T_1425 = $signed(io_boxYPosition_16) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1433 = $signed(io_boxXPosition_5) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_1434 = $signed(io_boxXPosition_17) < $signed(_T_73); // @[BoxDetection.scala 27:51]
  wire  _T_1435 = _T_1433 & _T_1434; // @[BoxDetection.scala 27:41]
  wire  _T_1436 = $signed(io_boxYPosition_5) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_1437 = _T_1435 & _T_1436; // @[BoxDetection.scala 27:60]
  wire  _T_1438 = $signed(io_boxYPosition_17) < $signed(_T_76); // @[BoxDetection.scala 28:35]
  wire  _T_1543 = $signed(io_boxXPosition_6) < $signed(_T_99); // @[BoxDetection.scala 27:32]
  wire  _T_1544 = $signed(io_boxXPosition_7) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1545 = _T_1543 & _T_1544; // @[BoxDetection.scala 27:41]
  wire  _T_1546 = $signed(io_boxYPosition_6) < $signed(_T_102); // @[BoxDetection.scala 28:16]
  wire  _T_1547 = _T_1545 & _T_1546; // @[BoxDetection.scala 27:60]
  wire  _T_1548 = $signed(io_boxYPosition_7) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1556 = $signed(io_boxXPosition_6) < $signed(_T_112); // @[BoxDetection.scala 27:32]
  wire  _T_1557 = $signed(io_boxXPosition_8) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1558 = _T_1556 & _T_1557; // @[BoxDetection.scala 27:41]
  wire  _T_1559 = $signed(io_boxYPosition_6) < $signed(_T_115); // @[BoxDetection.scala 28:16]
  wire  _T_1560 = _T_1558 & _T_1559; // @[BoxDetection.scala 27:60]
  wire  _T_1561 = $signed(io_boxYPosition_8) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1569 = $signed(io_boxXPosition_6) < $signed(_T_125); // @[BoxDetection.scala 27:32]
  wire  _T_1570 = $signed(io_boxXPosition_9) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1571 = _T_1569 & _T_1570; // @[BoxDetection.scala 27:41]
  wire  _T_1572 = $signed(io_boxYPosition_6) < $signed(_T_128); // @[BoxDetection.scala 28:16]
  wire  _T_1573 = _T_1571 & _T_1572; // @[BoxDetection.scala 27:60]
  wire  _T_1574 = $signed(io_boxYPosition_9) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1582 = $signed(io_boxXPosition_6) < $signed(_T_138); // @[BoxDetection.scala 27:32]
  wire  _T_1583 = $signed(io_boxXPosition_10) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1584 = _T_1582 & _T_1583; // @[BoxDetection.scala 27:41]
  wire  _T_1585 = $signed(io_boxYPosition_6) < $signed(_T_141); // @[BoxDetection.scala 28:16]
  wire  _T_1586 = _T_1584 & _T_1585; // @[BoxDetection.scala 27:60]
  wire  _T_1587 = $signed(io_boxYPosition_10) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1595 = $signed(io_boxXPosition_6) < $signed(_T_151); // @[BoxDetection.scala 27:32]
  wire  _T_1596 = $signed(io_boxXPosition_11) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1597 = _T_1595 & _T_1596; // @[BoxDetection.scala 27:41]
  wire  _T_1598 = $signed(io_boxYPosition_6) < $signed(_T_154); // @[BoxDetection.scala 28:16]
  wire  _T_1599 = _T_1597 & _T_1598; // @[BoxDetection.scala 27:60]
  wire  _T_1600 = $signed(io_boxYPosition_11) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1608 = $signed(io_boxXPosition_6) < $signed(_T_164); // @[BoxDetection.scala 27:32]
  wire  _T_1609 = $signed(io_boxXPosition_12) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1610 = _T_1608 & _T_1609; // @[BoxDetection.scala 27:41]
  wire  _T_1611 = $signed(io_boxYPosition_6) < $signed(_T_167); // @[BoxDetection.scala 28:16]
  wire  _T_1612 = _T_1610 & _T_1611; // @[BoxDetection.scala 27:60]
  wire  _T_1613 = $signed(io_boxYPosition_12) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1621 = $signed(io_boxXPosition_6) < $signed(_T_177); // @[BoxDetection.scala 27:32]
  wire  _T_1622 = $signed(io_boxXPosition_13) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1623 = _T_1621 & _T_1622; // @[BoxDetection.scala 27:41]
  wire  _T_1624 = $signed(io_boxYPosition_6) < $signed(_T_180); // @[BoxDetection.scala 28:16]
  wire  _T_1625 = _T_1623 & _T_1624; // @[BoxDetection.scala 27:60]
  wire  _T_1626 = $signed(io_boxYPosition_13) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1634 = $signed(io_boxXPosition_6) < $signed(_T_190); // @[BoxDetection.scala 27:32]
  wire  _T_1635 = $signed(io_boxXPosition_14) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1636 = _T_1634 & _T_1635; // @[BoxDetection.scala 27:41]
  wire  _T_1637 = $signed(io_boxYPosition_6) < $signed(_T_193); // @[BoxDetection.scala 28:16]
  wire  _T_1638 = _T_1636 & _T_1637; // @[BoxDetection.scala 27:60]
  wire  _T_1639 = $signed(io_boxYPosition_14) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1647 = $signed(io_boxXPosition_6) < $signed(_T_203); // @[BoxDetection.scala 27:32]
  wire  _T_1648 = $signed(io_boxXPosition_15) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1649 = _T_1647 & _T_1648; // @[BoxDetection.scala 27:41]
  wire  _T_1650 = $signed(io_boxYPosition_6) < $signed(_T_206); // @[BoxDetection.scala 28:16]
  wire  _T_1651 = _T_1649 & _T_1650; // @[BoxDetection.scala 27:60]
  wire  _T_1652 = $signed(io_boxYPosition_15) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  wire  _T_1673 = $signed(io_boxXPosition_6) < $signed(_T_229); // @[BoxDetection.scala 27:32]
  wire  _T_1674 = $signed(io_boxXPosition_17) < $signed(_T_86); // @[BoxDetection.scala 27:51]
  wire  _T_1675 = _T_1673 & _T_1674; // @[BoxDetection.scala 27:41]
  wire  _T_1676 = $signed(io_boxYPosition_6) < $signed(_T_232); // @[BoxDetection.scala 28:16]
  wire  _T_1677 = _T_1675 & _T_1676; // @[BoxDetection.scala 27:60]
  wire  _T_1678 = $signed(io_boxYPosition_17) < $signed(_T_89); // @[BoxDetection.scala 28:35]
  reg  _T_4320_0_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_0_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_2_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_3_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_4_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_16; // @[BoxDetection.scala 32:24]
  reg  _T_4320_5_17; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_7; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_8; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_9; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_10; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_11; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_12; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_13; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_14; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_15; // @[BoxDetection.scala 32:24]
  reg  _T_4320_6_17; // @[BoxDetection.scala 32:24]
  assign io_overlap_0_7 = _T_4320_0_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_8 = _T_4320_0_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_9 = _T_4320_0_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_10 = _T_4320_0_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_11 = _T_4320_0_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_12 = _T_4320_0_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_13 = _T_4320_0_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_14 = _T_4320_0_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_15 = _T_4320_0_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_16 = _T_4320_0_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_0_17 = _T_4320_0_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_7 = _T_4320_2_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_8 = _T_4320_2_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_9 = _T_4320_2_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_10 = _T_4320_2_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_11 = _T_4320_2_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_12 = _T_4320_2_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_13 = _T_4320_2_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_14 = _T_4320_2_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_15 = _T_4320_2_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_16 = _T_4320_2_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_2_17 = _T_4320_2_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_7 = _T_4320_3_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_8 = _T_4320_3_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_9 = _T_4320_3_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_10 = _T_4320_3_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_11 = _T_4320_3_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_12 = _T_4320_3_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_13 = _T_4320_3_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_14 = _T_4320_3_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_15 = _T_4320_3_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_16 = _T_4320_3_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_3_17 = _T_4320_3_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_7 = _T_4320_4_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_8 = _T_4320_4_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_9 = _T_4320_4_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_10 = _T_4320_4_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_11 = _T_4320_4_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_12 = _T_4320_4_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_13 = _T_4320_4_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_14 = _T_4320_4_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_15 = _T_4320_4_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_16 = _T_4320_4_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_4_17 = _T_4320_4_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_7 = _T_4320_5_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_8 = _T_4320_5_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_9 = _T_4320_5_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_10 = _T_4320_5_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_11 = _T_4320_5_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_12 = _T_4320_5_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_13 = _T_4320_5_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_14 = _T_4320_5_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_15 = _T_4320_5_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_16 = _T_4320_5_16; // @[BoxDetection.scala 32:14]
  assign io_overlap_5_17 = _T_4320_5_17; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_7 = _T_4320_6_7; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_8 = _T_4320_6_8; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_9 = _T_4320_6_9; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_10 = _T_4320_6_10; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_11 = _T_4320_6_11; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_12 = _T_4320_6_12; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_13 = _T_4320_6_13; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_14 = _T_4320_6_14; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_15 = _T_4320_6_15; // @[BoxDetection.scala 32:14]
  assign io_overlap_6_17 = _T_4320_6_17; // @[BoxDetection.scala 32:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4320_0_7 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_4320_0_8 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_4320_0_9 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_4320_0_10 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_4320_0_11 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_4320_0_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_4320_0_13 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_4320_0_14 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_4320_0_15 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_4320_0_16 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_4320_0_17 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_4320_2_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_4320_2_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_4320_2_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_4320_2_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_4320_2_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_4320_2_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_4320_2_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_4320_2_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_4320_2_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_4320_2_16 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4320_2_17 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4320_3_7 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4320_3_8 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4320_3_9 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4320_3_10 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4320_3_11 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4320_3_12 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4320_3_13 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4320_3_14 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4320_3_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4320_3_16 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4320_3_17 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4320_4_7 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4320_4_8 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4320_4_9 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4320_4_10 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4320_4_11 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4320_4_12 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4320_4_13 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4320_4_14 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4320_4_15 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4320_4_16 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4320_4_17 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4320_5_7 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4320_5_8 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4320_5_9 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4320_5_10 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4320_5_11 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4320_5_12 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4320_5_13 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4320_5_14 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4320_5_15 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4320_5_16 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4320_5_17 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4320_6_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4320_6_8 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4320_6_9 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4320_6_10 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4320_6_11 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4320_6_12 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4320_6_13 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4320_6_14 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4320_6_15 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4320_6_17 = _RAND_64[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_4320_0_7 <= _T_107 & _T_108;
    _T_4320_0_8 <= _T_120 & _T_121;
    _T_4320_0_9 <= _T_133 & _T_134;
    _T_4320_0_10 <= _T_146 & _T_147;
    _T_4320_0_11 <= _T_159 & _T_160;
    _T_4320_0_12 <= _T_172 & _T_173;
    _T_4320_0_13 <= _T_185 & _T_186;
    _T_4320_0_14 <= _T_198 & _T_199;
    _T_4320_0_15 <= _T_211 & _T_212;
    _T_4320_0_16 <= _T_224 & _T_225;
    _T_4320_0_17 <= _T_237 & _T_238;
    _T_4320_2_7 <= _T_587 & _T_588;
    _T_4320_2_8 <= _T_600 & _T_601;
    _T_4320_2_9 <= _T_613 & _T_614;
    _T_4320_2_10 <= _T_626 & _T_627;
    _T_4320_2_11 <= _T_639 & _T_640;
    _T_4320_2_12 <= _T_652 & _T_653;
    _T_4320_2_13 <= _T_665 & _T_666;
    _T_4320_2_14 <= _T_678 & _T_679;
    _T_4320_2_15 <= _T_691 & _T_692;
    _T_4320_2_16 <= _T_704 & _T_705;
    _T_4320_2_17 <= _T_717 & _T_718;
    _T_4320_3_7 <= _T_827 & _T_828;
    _T_4320_3_8 <= _T_840 & _T_841;
    _T_4320_3_9 <= _T_853 & _T_854;
    _T_4320_3_10 <= _T_866 & _T_867;
    _T_4320_3_11 <= _T_879 & _T_880;
    _T_4320_3_12 <= _T_892 & _T_893;
    _T_4320_3_13 <= _T_905 & _T_906;
    _T_4320_3_14 <= _T_918 & _T_919;
    _T_4320_3_15 <= _T_931 & _T_932;
    _T_4320_3_16 <= _T_944 & _T_945;
    _T_4320_3_17 <= _T_957 & _T_958;
    _T_4320_4_7 <= _T_1067 & _T_1068;
    _T_4320_4_8 <= _T_1080 & _T_1081;
    _T_4320_4_9 <= _T_1093 & _T_1094;
    _T_4320_4_10 <= _T_1106 & _T_1107;
    _T_4320_4_11 <= _T_1119 & _T_1120;
    _T_4320_4_12 <= _T_1132 & _T_1133;
    _T_4320_4_13 <= _T_1145 & _T_1146;
    _T_4320_4_14 <= _T_1158 & _T_1159;
    _T_4320_4_15 <= _T_1171 & _T_1172;
    _T_4320_4_16 <= _T_1184 & _T_1185;
    _T_4320_4_17 <= _T_1197 & _T_1198;
    _T_4320_5_7 <= _T_1307 & _T_1308;
    _T_4320_5_8 <= _T_1320 & _T_1321;
    _T_4320_5_9 <= _T_1333 & _T_1334;
    _T_4320_5_10 <= _T_1346 & _T_1347;
    _T_4320_5_11 <= _T_1359 & _T_1360;
    _T_4320_5_12 <= _T_1372 & _T_1373;
    _T_4320_5_13 <= _T_1385 & _T_1386;
    _T_4320_5_14 <= _T_1398 & _T_1399;
    _T_4320_5_15 <= _T_1411 & _T_1412;
    _T_4320_5_16 <= _T_1424 & _T_1425;
    _T_4320_5_17 <= _T_1437 & _T_1438;
    _T_4320_6_7 <= _T_1547 & _T_1548;
    _T_4320_6_8 <= _T_1560 & _T_1561;
    _T_4320_6_9 <= _T_1573 & _T_1574;
    _T_4320_6_10 <= _T_1586 & _T_1587;
    _T_4320_6_11 <= _T_1599 & _T_1600;
    _T_4320_6_12 <= _T_1612 & _T_1613;
    _T_4320_6_13 <= _T_1625 & _T_1626;
    _T_4320_6_14 <= _T_1638 & _T_1639;
    _T_4320_6_15 <= _T_1651 & _T_1652;
    _T_4320_6_17 <= _T_1677 & _T_1678;
  end
endmodule
module Randomizer(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_1(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_2(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h8;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_3(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h8;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_4(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h9;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_5(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h9;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_6(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'ha;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_7(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'ha;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_8(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hb;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_9(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hb;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_10(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hc;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_11(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hc;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_12(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hd;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_13(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hd;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_14(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'he;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_15(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'he;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_16(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hf;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_17(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'hf;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_18(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h10;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_19(
  input        clock,
  input        reset,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [6:0] place; // @[Randomizer.scala 19:22]
  reg [6:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 7'h40; // @[Randomizer.scala 26:14]
  wire [7:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h10;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 7'h0;
    end else begin
      place <= {{1'd0}, state[5:0]};
    end
    if (reset) begin
      placeholder <= 7'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[6:0];
    end
  end
endmodule
module Randomizer_33(
  input        clock,
  input        reset,
  output [1:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [1:0] place; // @[Randomizer.scala 19:22]
  reg [1:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 2'h2; // @[Randomizer.scala 26:14]
  wire [2:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h1;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 2'h0;
    end else begin
      place <= {{1'd0}, state[0]};
    end
    if (reset) begin
      placeholder <= 2'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[1:0];
    end
  end
endmodule
module Randomizer_34(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7d;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_35(
  input        clock,
  input        reset,
  output [5:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [5:0] place; // @[Randomizer.scala 19:22]
  reg [5:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 6'h11; // @[Randomizer.scala 26:14]
  wire [6:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h9;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 6'h0;
    end else begin
      place <= {{1'd0}, state[4:0]};
    end
    if (reset) begin
      placeholder <= 6'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[5:0];
    end
  end
endmodule
module Randomizer_36(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7e;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_38(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7f;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_40(
  input        clock,
  input        reset,
  output [1:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [1:0] place; // @[Randomizer.scala 19:22]
  reg [1:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 2'h2; // @[Randomizer.scala 26:14]
  wire [2:0] _T_14 = {{1'd0}, place}; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h2;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 2'h0;
    end else begin
      place <= {{1'd0}, state[0]};
    end
    if (reset) begin
      placeholder <= 2'h0;
    end else if (_T_11) begin
      placeholder <= _T_14[1:0];
    end
  end
endmodule
module Randomizer_41(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7a;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_43(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7b;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module Randomizer_45(
  input        clock,
  input        reset,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] state; // @[Randomizer.scala 13:22]
  wire [8:0] _T_1 = {{4'd0}, state[8:4]}; // @[Randomizer.scala 16:32]
  wire [8:0] _T_2 = state ^ _T_1; // @[Randomizer.scala 16:23]
  wire [8:0] _T_3 = {{5'd0}, state[8:5]}; // @[Randomizer.scala 16:49]
  wire [8:0] _T_4 = _T_2 ^ _T_3; // @[Randomizer.scala 16:40]
  wire [8:0] _T_5 = {{6'd0}, state[8:6]}; // @[Randomizer.scala 16:66]
  wire [8:0] _T_6 = _T_4 ^ _T_5; // @[Randomizer.scala 16:57]
  wire [8:0] newbit = _T_6 & 9'h1; // @[Randomizer.scala 16:75]
  wire [8:0] _T_7 = {{1'd0}, state[8:1]}; // @[Randomizer.scala 17:19]
  wire [16:0] _GEN_5 = {newbit, 8'h0}; // @[Randomizer.scala 17:37]
  wire [23:0] _T_8 = {{7'd0}, _GEN_5}; // @[Randomizer.scala 17:37]
  wire [23:0] _GEN_6 = {{15'd0}, _T_7}; // @[Randomizer.scala 17:27]
  wire [23:0] _T_9 = _GEN_6 | _T_8; // @[Randomizer.scala 17:27]
  reg [9:0] place; // @[Randomizer.scala 19:22]
  reg [9:0] placeholder; // @[Randomizer.scala 21:28]
  wire  _T_11 = place <= 10'h100; // @[Randomizer.scala 26:14]
  wire [9:0] _T_15 = place + 10'h60; // @[Randomizer.scala 27:26]
  assign io_out = placeholder; // @[Randomizer.scala 30:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  place = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  placeholder = _RAND_2[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 9'h7c;
    end else begin
      state <= _T_9[8:0];
    end
    if (reset) begin
      place <= 10'h0;
    end else begin
      place <= {{2'd0}, state[7:0]};
    end
    if (reset) begin
      placeholder <= 10'h0;
    end else if (_T_11) begin
      placeholder <= _T_15;
    end
  end
endmodule
module GameLogic(
  input         clock,
  input         reset,
  input         io_btnC,
  input         io_btnU,
  input         io_btnL,
  input         io_btnR,
  input         io_btnD,
  input         io_sw_0,
  input         io_sw_1,
  input         io_sw_2,
  input         io_sw_7,
  output [3:0]  io_songInput,
  output [10:0] io_spriteXPosition_0,
  output [10:0] io_spriteXPosition_1,
  output [10:0] io_spriteXPosition_2,
  output [10:0] io_spriteXPosition_3,
  output [10:0] io_spriteXPosition_4,
  output [10:0] io_spriteXPosition_5,
  output [10:0] io_spriteXPosition_6,
  output [10:0] io_spriteXPosition_7,
  output [10:0] io_spriteXPosition_8,
  output [10:0] io_spriteXPosition_9,
  output [10:0] io_spriteXPosition_10,
  output [10:0] io_spriteXPosition_11,
  output [10:0] io_spriteXPosition_12,
  output [10:0] io_spriteXPosition_13,
  output [10:0] io_spriteXPosition_14,
  output [10:0] io_spriteXPosition_15,
  output [10:0] io_spriteXPosition_16,
  output [10:0] io_spriteXPosition_17,
  output [10:0] io_spriteXPosition_18,
  output [10:0] io_spriteXPosition_19,
  output [10:0] io_spriteXPosition_20,
  output [10:0] io_spriteXPosition_21,
  output [10:0] io_spriteXPosition_22,
  output [10:0] io_spriteXPosition_23,
  output [10:0] io_spriteXPosition_24,
  output [10:0] io_spriteXPosition_25,
  output [10:0] io_spriteXPosition_26,
  output [10:0] io_spriteXPosition_27,
  output [10:0] io_spriteXPosition_28,
  output [10:0] io_spriteXPosition_29,
  output [10:0] io_spriteXPosition_30,
  output [10:0] io_spriteXPosition_31,
  output [10:0] io_spriteXPosition_32,
  output [10:0] io_spriteXPosition_33,
  output [10:0] io_spriteXPosition_41,
  output [10:0] io_spriteXPosition_42,
  output [10:0] io_spriteXPosition_43,
  output [10:0] io_spriteXPosition_44,
  output [10:0] io_spriteXPosition_45,
  output [10:0] io_spriteXPosition_46,
  output [10:0] io_spriteXPosition_47,
  output [10:0] io_spriteXPosition_48,
  output [10:0] io_spriteXPosition_49,
  output [10:0] io_spriteXPosition_50,
  output [10:0] io_spriteXPosition_51,
  output [10:0] io_spriteXPosition_122,
  output [10:0] io_spriteXPosition_123,
  output [10:0] io_spriteXPosition_124,
  output [10:0] io_spriteXPosition_125,
  output [10:0] io_spriteXPosition_126,
  output [10:0] io_spriteXPosition_127,
  output [9:0]  io_spriteYPosition_0,
  output [9:0]  io_spriteYPosition_1,
  output [9:0]  io_spriteYPosition_2,
  output [9:0]  io_spriteYPosition_3,
  output [9:0]  io_spriteYPosition_4,
  output [9:0]  io_spriteYPosition_5,
  output [9:0]  io_spriteYPosition_6,
  output [9:0]  io_spriteYPosition_7,
  output [9:0]  io_spriteYPosition_8,
  output [9:0]  io_spriteYPosition_9,
  output [9:0]  io_spriteYPosition_10,
  output [9:0]  io_spriteYPosition_11,
  output [9:0]  io_spriteYPosition_12,
  output [9:0]  io_spriteYPosition_13,
  output [9:0]  io_spriteYPosition_14,
  output [9:0]  io_spriteYPosition_15,
  output [9:0]  io_spriteYPosition_16,
  output [9:0]  io_spriteYPosition_17,
  output [9:0]  io_spriteYPosition_18,
  output [9:0]  io_spriteYPosition_19,
  output [9:0]  io_spriteYPosition_20,
  output [9:0]  io_spriteYPosition_21,
  output [9:0]  io_spriteYPosition_22,
  output [9:0]  io_spriteYPosition_23,
  output [9:0]  io_spriteYPosition_24,
  output [9:0]  io_spriteYPosition_25,
  output [9:0]  io_spriteYPosition_26,
  output [9:0]  io_spriteYPosition_27,
  output [9:0]  io_spriteYPosition_28,
  output [9:0]  io_spriteYPosition_29,
  output [9:0]  io_spriteYPosition_30,
  output [9:0]  io_spriteYPosition_31,
  output [9:0]  io_spriteYPosition_32,
  output [9:0]  io_spriteYPosition_33,
  output [9:0]  io_spriteYPosition_41,
  output [9:0]  io_spriteYPosition_42,
  output [9:0]  io_spriteYPosition_43,
  output [9:0]  io_spriteYPosition_122,
  output [9:0]  io_spriteYPosition_123,
  output [9:0]  io_spriteYPosition_124,
  output [9:0]  io_spriteYPosition_125,
  output [9:0]  io_spriteYPosition_126,
  output [9:0]  io_spriteYPosition_127,
  output        io_spriteVisible_0,
  output        io_spriteVisible_1,
  output        io_spriteVisible_2,
  output        io_spriteVisible_3,
  output        io_spriteVisible_4,
  output        io_spriteVisible_5,
  output        io_spriteVisible_6,
  output        io_spriteVisible_7,
  output        io_spriteVisible_8,
  output        io_spriteVisible_9,
  output        io_spriteVisible_10,
  output        io_spriteVisible_11,
  output        io_spriteVisible_12,
  output        io_spriteVisible_13,
  output        io_spriteVisible_14,
  output        io_spriteVisible_15,
  output        io_spriteVisible_16,
  output        io_spriteVisible_17,
  output        io_spriteVisible_18,
  output        io_spriteVisible_19,
  output        io_spriteVisible_20,
  output        io_spriteVisible_21,
  output        io_spriteVisible_22,
  output        io_spriteVisible_23,
  output        io_spriteVisible_24,
  output        io_spriteVisible_25,
  output        io_spriteVisible_26,
  output        io_spriteVisible_27,
  output        io_spriteVisible_28,
  output        io_spriteVisible_29,
  output        io_spriteVisible_30,
  output        io_spriteVisible_31,
  output        io_spriteVisible_32,
  output        io_spriteVisible_33,
  output        io_spriteVisible_41,
  output        io_spriteVisible_42,
  output        io_spriteVisible_43,
  output        io_spriteVisible_44,
  output        io_spriteVisible_45,
  output        io_spriteVisible_46,
  output        io_spriteVisible_47,
  output        io_spriteVisible_48,
  output        io_spriteVisible_49,
  output        io_spriteVisible_50,
  output        io_spriteVisible_51,
  output        io_spriteVisible_55,
  output        io_spriteVisible_56,
  output        io_spriteVisible_57,
  output        io_spriteVisible_61,
  output        io_spriteVisible_62,
  output        io_spriteVisible_63,
  output        io_spriteVisible_64,
  output        io_spriteVisible_65,
  output        io_spriteVisible_66,
  output        io_spriteVisible_70,
  output        io_spriteVisible_71,
  output        io_spriteVisible_72,
  output        io_spriteFlipVertical_122,
  output        io_spriteFlipVertical_123,
  output        io_spriteFlipVertical_124,
  output        io_spriteFlipVertical_125,
  output        io_spriteFlipVertical_126,
  output        io_spriteFlipVertical_127,
  output [9:0]  io_viewBoxX_0,
  output [4:0]  io_backBufferWriteData,
  output [10:0] io_backBufferWriteAddress,
  output        io_backBufferWriteEnable,
  input         io_newFrame,
  output        io_frameUpdateDone
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
`endif // RANDOMIZE_REG_INIT
  wire  boxDetection_clock; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_0; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_2; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_3; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_4; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_5; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_6; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_7; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_8; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_9; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_10; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_11; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_12; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_13; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_14; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_15; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_16; // @[GameLogic.scala 700:28]
  wire [10:0] boxDetection_io_boxXPosition_17; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_0; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_2; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_3; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_4; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_5; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_6; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_7; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_8; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_9; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_10; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_11; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_12; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_13; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_14; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_15; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_16; // @[GameLogic.scala 700:28]
  wire [9:0] boxDetection_io_boxYPosition_17; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_7; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_8; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_9; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_10; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_11; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_12; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_13; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_14; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_15; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_16; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_0_17; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_7; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_8; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_9; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_10; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_11; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_12; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_13; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_14; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_15; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_16; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_2_17; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_7; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_8; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_9; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_10; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_11; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_12; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_13; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_14; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_15; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_16; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_3_17; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_7; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_8; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_9; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_10; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_11; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_12; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_13; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_14; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_15; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_16; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_4_17; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_7; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_8; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_9; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_10; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_11; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_12; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_13; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_14; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_15; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_16; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_5_17; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_7; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_8; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_9; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_10; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_11; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_12; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_13; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_14; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_15; // @[GameLogic.scala 700:28]
  wire  boxDetection_io_overlap_6_17; // @[GameLogic.scala 700:28]
  wire  Randomizer_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_1_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_1_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_1_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_2_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_2_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_2_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_3_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_3_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_3_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_4_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_4_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_4_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_5_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_5_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_5_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_6_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_6_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_6_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_7_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_7_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_7_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_8_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_8_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_8_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_9_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_9_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_9_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_10_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_10_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_10_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_11_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_11_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_11_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_12_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_12_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_12_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_13_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_13_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_13_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_14_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_14_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_14_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_15_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_15_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_15_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_16_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_16_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_16_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_17_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_17_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_17_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_18_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_18_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_18_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_19_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_19_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_19_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_20_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_20_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_20_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_21_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_21_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_21_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_22_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_22_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_22_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_23_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_23_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_23_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_24_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_24_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_24_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_25_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_25_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_25_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_26_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_26_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_26_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_27_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_27_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_27_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_28_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_28_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_28_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_29_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_29_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_29_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_30_clock; // @[GameLogic.scala 189:24]
  wire  Randomizer_30_reset; // @[GameLogic.scala 189:24]
  wire [9:0] Randomizer_30_io_out; // @[GameLogic.scala 189:24]
  wire  Randomizer_31_clock; // @[GameLogic.scala 190:31]
  wire  Randomizer_31_reset; // @[GameLogic.scala 190:31]
  wire [6:0] Randomizer_31_io_out; // @[GameLogic.scala 190:31]
  wire  Randomizer_32_clock; // @[GameLogic.scala 362:24]
  wire  Randomizer_32_reset; // @[GameLogic.scala 362:24]
  wire [9:0] Randomizer_32_io_out; // @[GameLogic.scala 362:24]
  wire  Randomizer_33_clock; // @[GameLogic.scala 118:24]
  wire  Randomizer_33_reset; // @[GameLogic.scala 118:24]
  wire [1:0] Randomizer_33_io_out; // @[GameLogic.scala 118:24]
  wire  Randomizer_34_clock; // @[GameLogic.scala 95:24]
  wire  Randomizer_34_reset; // @[GameLogic.scala 95:24]
  wire [9:0] Randomizer_34_io_out; // @[GameLogic.scala 95:24]
  wire  Randomizer_35_clock; // @[GameLogic.scala 96:25]
  wire  Randomizer_35_reset; // @[GameLogic.scala 96:25]
  wire [5:0] Randomizer_35_io_out; // @[GameLogic.scala 96:25]
  wire  Randomizer_36_clock; // @[GameLogic.scala 95:24]
  wire  Randomizer_36_reset; // @[GameLogic.scala 95:24]
  wire [9:0] Randomizer_36_io_out; // @[GameLogic.scala 95:24]
  wire  Randomizer_37_clock; // @[GameLogic.scala 96:25]
  wire  Randomizer_37_reset; // @[GameLogic.scala 96:25]
  wire [5:0] Randomizer_37_io_out; // @[GameLogic.scala 96:25]
  wire  Randomizer_38_clock; // @[GameLogic.scala 95:24]
  wire  Randomizer_38_reset; // @[GameLogic.scala 95:24]
  wire [9:0] Randomizer_38_io_out; // @[GameLogic.scala 95:24]
  wire  Randomizer_39_clock; // @[GameLogic.scala 96:25]
  wire  Randomizer_39_reset; // @[GameLogic.scala 96:25]
  wire [5:0] Randomizer_39_io_out; // @[GameLogic.scala 96:25]
  wire  Randomizer_40_clock; // @[GameLogic.scala 118:24]
  wire  Randomizer_40_reset; // @[GameLogic.scala 118:24]
  wire [1:0] Randomizer_40_io_out; // @[GameLogic.scala 118:24]
  wire  Randomizer_41_clock; // @[GameLogic.scala 95:24]
  wire  Randomizer_41_reset; // @[GameLogic.scala 95:24]
  wire [9:0] Randomizer_41_io_out; // @[GameLogic.scala 95:24]
  wire  Randomizer_42_clock; // @[GameLogic.scala 96:25]
  wire  Randomizer_42_reset; // @[GameLogic.scala 96:25]
  wire [5:0] Randomizer_42_io_out; // @[GameLogic.scala 96:25]
  wire  Randomizer_43_clock; // @[GameLogic.scala 95:24]
  wire  Randomizer_43_reset; // @[GameLogic.scala 95:24]
  wire [9:0] Randomizer_43_io_out; // @[GameLogic.scala 95:24]
  wire  Randomizer_44_clock; // @[GameLogic.scala 96:25]
  wire  Randomizer_44_reset; // @[GameLogic.scala 96:25]
  wire [5:0] Randomizer_44_io_out; // @[GameLogic.scala 96:25]
  wire  Randomizer_45_clock; // @[GameLogic.scala 95:24]
  wire  Randomizer_45_reset; // @[GameLogic.scala 95:24]
  wire [9:0] Randomizer_45_io_out; // @[GameLogic.scala 95:24]
  wire  Randomizer_46_clock; // @[GameLogic.scala 96:25]
  wire  Randomizer_46_reset; // @[GameLogic.scala 96:25]
  wire [5:0] Randomizer_46_io_out; // @[GameLogic.scala 96:25]
  reg  planetUp; // @[GameLogic.scala 347:25]
  reg [10:0] Xstart_0; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_1; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_2; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_3; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_4; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_5; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_6; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_7; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_8; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_9; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_10; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_11; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_12; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_13; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_14; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_15; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_16; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_17; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_18; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_19; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_20; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_21; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_22; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_23; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_24; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_25; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_26; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_27; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_28; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_29; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_30; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_31; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_32; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_33; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_41; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_42; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_43; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_44; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_45; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_46; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_47; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_48; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_49; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_50; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_51; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_122; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_123; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_124; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_125; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_126; // @[GameLogic.scala 412:23]
  reg [10:0] Xstart_127; // @[GameLogic.scala 412:23]
  reg [10:0] Ystart_0; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_1; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_2; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_3; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_4; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_5; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_6; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_7; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_8; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_9; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_10; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_11; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_12; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_13; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_14; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_15; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_16; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_17; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_18; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_19; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_20; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_21; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_22; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_23; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_24; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_25; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_26; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_27; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_28; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_29; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_30; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_31; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_32; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_33; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_41; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_42; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_43; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_122; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_123; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_124; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_125; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_126; // @[GameLogic.scala 497:23]
  reg [10:0] Ystart_127; // @[GameLogic.scala 497:23]
  reg  spriteVisibleReg_0; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_1; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_2; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_3; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_4; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_5; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_6; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_7; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_8; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_9; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_10; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_11; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_12; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_13; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_14; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_15; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_16; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_17; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_18; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_19; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_20; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_21; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_22; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_23; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_24; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_25; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_26; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_27; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_28; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_29; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_30; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_31; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_32; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_33; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_41; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_42; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_43; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_44; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_45; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_46; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_47; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_48; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_49; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_50; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_51; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_55; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_56; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_57; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_61; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_62; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_63; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_64; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_65; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_66; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_70; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_71; // @[GameLogic.scala 608:33]
  reg  spriteVisibleReg_72; // @[GameLogic.scala 608:33]
  reg  spriteFlipVerticalReg_122; // @[GameLogic.scala 610:38]
  reg  spriteFlipVerticalReg_123; // @[GameLogic.scala 610:38]
  reg  spriteFlipVerticalReg_124; // @[GameLogic.scala 610:38]
  reg  spriteFlipVerticalReg_125; // @[GameLogic.scala 610:38]
  reg  spriteFlipVerticalReg_126; // @[GameLogic.scala 610:38]
  reg  spriteFlipVerticalReg_127; // @[GameLogic.scala 610:38]
  reg  btnCReg; // @[GameLogic.scala 611:24]
  reg [9:0] viewX; // @[GameLogic.scala 636:22]
  reg [3:0] stateReg; // @[GameLogic.scala 655:25]
  reg [9:0] shotCnt; // @[GameLogic.scala 658:24]
  reg  shotLoad; // @[GameLogic.scala 659:25]
  reg [2:0] shotCntBig; // @[GameLogic.scala 660:27]
  reg [2:0] shotCntFast; // @[GameLogic.scala 661:28]
  reg  shotPop_0; // @[GameLogic.scala 662:24]
  reg  shotPop_1; // @[GameLogic.scala 662:24]
  reg  shotPop_2; // @[GameLogic.scala 662:24]
  reg  shotPop_3; // @[GameLogic.scala 662:24]
  reg  shotPop_4; // @[GameLogic.scala 662:24]
  reg  shotInteract_0; // @[GameLogic.scala 663:29]
  reg  shotInteract_1; // @[GameLogic.scala 663:29]
  reg  shotInteract_2; // @[GameLogic.scala 663:29]
  reg  shotInteract_3; // @[GameLogic.scala 663:29]
  reg  shotInteract_4; // @[GameLogic.scala 663:29]
  reg  astInteract_0; // @[GameLogic.scala 664:28]
  reg  astInteract_1; // @[GameLogic.scala 664:28]
  reg  astInteract_2; // @[GameLogic.scala 664:28]
  reg  astInteract_3; // @[GameLogic.scala 664:28]
  reg  astInteract_4; // @[GameLogic.scala 664:28]
  reg  astInteract_5; // @[GameLogic.scala 664:28]
  reg  astInteract_6; // @[GameLogic.scala 664:28]
  reg  astInteract_7; // @[GameLogic.scala 664:28]
  reg  astInteract_8; // @[GameLogic.scala 664:28]
  reg  astInteract_9; // @[GameLogic.scala 664:28]
  reg  astInteract_10; // @[GameLogic.scala 664:28]
  reg  shipInteract; // @[GameLogic.scala 665:29]
  reg  die_0; // @[GameLogic.scala 667:20]
  reg  die_1; // @[GameLogic.scala 667:20]
  reg  die_2; // @[GameLogic.scala 667:20]
  reg  die_3; // @[GameLogic.scala 667:20]
  reg  die_4; // @[GameLogic.scala 667:20]
  reg  die_5; // @[GameLogic.scala 667:20]
  reg  die_6; // @[GameLogic.scala 667:20]
  reg  die_7; // @[GameLogic.scala 667:20]
  reg  die_8; // @[GameLogic.scala 667:20]
  reg  die_9; // @[GameLogic.scala 667:20]
  reg  die_10; // @[GameLogic.scala 667:20]
  reg  kill_0_0; // @[GameLogic.scala 668:21]
  reg  kill_0_1; // @[GameLogic.scala 668:21]
  reg  kill_0_2; // @[GameLogic.scala 668:21]
  reg  kill_0_3; // @[GameLogic.scala 668:21]
  reg  kill_0_4; // @[GameLogic.scala 668:21]
  reg  kill_1_0; // @[GameLogic.scala 668:21]
  reg  kill_1_1; // @[GameLogic.scala 668:21]
  reg  kill_1_2; // @[GameLogic.scala 668:21]
  reg  kill_1_3; // @[GameLogic.scala 668:21]
  reg  kill_1_4; // @[GameLogic.scala 668:21]
  reg  kill_2_0; // @[GameLogic.scala 668:21]
  reg  kill_2_1; // @[GameLogic.scala 668:21]
  reg  kill_2_2; // @[GameLogic.scala 668:21]
  reg  kill_2_3; // @[GameLogic.scala 668:21]
  reg  kill_2_4; // @[GameLogic.scala 668:21]
  reg  kill_3_0; // @[GameLogic.scala 668:21]
  reg  kill_3_1; // @[GameLogic.scala 668:21]
  reg  kill_3_2; // @[GameLogic.scala 668:21]
  reg  kill_3_3; // @[GameLogic.scala 668:21]
  reg  kill_3_4; // @[GameLogic.scala 668:21]
  reg  kill_4_0; // @[GameLogic.scala 668:21]
  reg  kill_4_1; // @[GameLogic.scala 668:21]
  reg  kill_4_2; // @[GameLogic.scala 668:21]
  reg  kill_4_3; // @[GameLogic.scala 668:21]
  reg  kill_4_4; // @[GameLogic.scala 668:21]
  reg  kill_5_0; // @[GameLogic.scala 668:21]
  reg  kill_5_1; // @[GameLogic.scala 668:21]
  reg  kill_5_2; // @[GameLogic.scala 668:21]
  reg  kill_5_3; // @[GameLogic.scala 668:21]
  reg  kill_5_4; // @[GameLogic.scala 668:21]
  reg  kill_6_0; // @[GameLogic.scala 668:21]
  reg  kill_6_1; // @[GameLogic.scala 668:21]
  reg  kill_6_2; // @[GameLogic.scala 668:21]
  reg  kill_6_3; // @[GameLogic.scala 668:21]
  reg  kill_6_4; // @[GameLogic.scala 668:21]
  reg  kill_7_0; // @[GameLogic.scala 668:21]
  reg  kill_7_1; // @[GameLogic.scala 668:21]
  reg  kill_7_2; // @[GameLogic.scala 668:21]
  reg  kill_7_3; // @[GameLogic.scala 668:21]
  reg  kill_7_4; // @[GameLogic.scala 668:21]
  reg  kill_8_0; // @[GameLogic.scala 668:21]
  reg  kill_8_1; // @[GameLogic.scala 668:21]
  reg  kill_8_2; // @[GameLogic.scala 668:21]
  reg  kill_8_3; // @[GameLogic.scala 668:21]
  reg  kill_8_4; // @[GameLogic.scala 668:21]
  reg  kill_9_0; // @[GameLogic.scala 668:21]
  reg  kill_9_1; // @[GameLogic.scala 668:21]
  reg  kill_9_2; // @[GameLogic.scala 668:21]
  reg  kill_9_3; // @[GameLogic.scala 668:21]
  reg  kill_10_0; // @[GameLogic.scala 668:21]
  reg  kill_10_1; // @[GameLogic.scala 668:21]
  reg  kill_10_2; // @[GameLogic.scala 668:21]
  reg  kill_10_3; // @[GameLogic.scala 668:21]
  reg  kill_10_4; // @[GameLogic.scala 668:21]
  reg [3:0] hp; // @[GameLogic.scala 670:19]
  reg [4:0] planetHp; // @[GameLogic.scala 671:25]
  reg [5:0] spwnProt; // @[GameLogic.scala 672:25]
  reg  show; // @[GameLogic.scala 673:21]
  reg  blink; // @[GameLogic.scala 674:22]
  reg [7:0] secCnt; // @[GameLogic.scala 675:23]
  reg [2:0] level; // @[GameLogic.scala 676:22]
  reg  start; // @[GameLogic.scala 677:22]
  reg  levelCng; // @[GameLogic.scala 678:25]
  reg [3:0] cngCnt; // @[GameLogic.scala 679:23]
  reg [9:0] cnt; // @[GameLogic.scala 681:20]
  wire  _T_24 = $signed(cnt) == 10'sh1d; // @[GameLogic.scala 682:17]
  wire  _T_25 = $signed(cnt) == 10'sh3b; // @[GameLogic.scala 682:33]
  wire  cng = _T_24 | _T_25; // @[GameLogic.scala 682:26]
  reg [6:0] count1; // @[GameLogic.scala 686:23]
  reg [6:0] count3; // @[GameLogic.scala 688:23]
  reg [7:0] count4; // @[GameLogic.scala 689:23]
  reg [7:0] count5; // @[GameLogic.scala 690:23]
  wire  _T_26 = ~show; // @[GameLogic.scala 694:26]
  wire  _T_27 = ~shipInteract; // @[GameLogic.scala 696:8]
  wire  _T_28 = _T_27 & blink; // @[GameLogic.scala 696:22]
  wire  _GEN_0 = _T_28 ? 1'h0 : show; // @[GameLogic.scala 696:32]
  wire  _GEN_1 = _T_28 ? 1'h0 : _T_26; // @[GameLogic.scala 696:32]
  wire [8:0] _T_32 = 8'sh0 / 8'sh2; // @[GameLogic.scala 702:66]
  wire [10:0] _GEN_4379 = {{2{_T_32[8]}},_T_32}; // @[GameLogic.scala 702:51]
  wire [10:0] _T_42 = $signed(Ystart_0) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_70 = $signed(Ystart_2) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_84 = $signed(Ystart_3) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_98 = $signed(Ystart_4) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_112 = $signed(Ystart_5) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_126 = $signed(Ystart_6) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [7:0] _T_129 = 8'sh20 - 8'sh8; // @[GameLogic.scala 702:57]
  wire [8:0] _T_130 = $signed(_T_129) / 8'sh2; // @[GameLogic.scala 702:66]
  wire [10:0] _GEN_4393 = {{2{_T_130[8]}},_T_130}; // @[GameLogic.scala 702:51]
  wire [10:0] _T_140 = $signed(Ystart_7) + $signed(_GEN_4393); // @[GameLogic.scala 703:51]
  wire [7:0] _T_143 = 8'sh20 - 8'sh10; // @[GameLogic.scala 702:57]
  wire [8:0] _T_144 = $signed(_T_143) / 8'sh2; // @[GameLogic.scala 702:66]
  wire [10:0] _GEN_4395 = {{2{_T_144[8]}},_T_144}; // @[GameLogic.scala 702:51]
  wire [10:0] _T_154 = $signed(Ystart_8) + $signed(_GEN_4395); // @[GameLogic.scala 703:51]
  wire [7:0] _T_157 = 8'sh20 - 8'sh1c; // @[GameLogic.scala 702:57]
  wire [8:0] _T_158 = $signed(_T_157) / 8'sh2; // @[GameLogic.scala 702:66]
  wire [10:0] _GEN_4397 = {{2{_T_158[8]}},_T_158}; // @[GameLogic.scala 702:51]
  wire [10:0] _T_168 = $signed(Ystart_9) + $signed(_GEN_4397); // @[GameLogic.scala 703:51]
  wire [10:0] _T_182 = $signed(Ystart_10) + $signed(_GEN_4397); // @[GameLogic.scala 703:51]
  wire [10:0] _T_196 = $signed(Ystart_11) + $signed(_GEN_4397); // @[GameLogic.scala 703:51]
  wire [10:0] _T_210 = $signed(Ystart_12) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_224 = $signed(Ystart_13) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_238 = $signed(Ystart_14) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_252 = $signed(Ystart_15) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [10:0] _T_266 = $signed(Ystart_16) + $signed(_GEN_4379); // @[GameLogic.scala 703:51]
  wire [7:0] _T_269 = 8'sh20 - 8'sh60; // @[GameLogic.scala 702:57]
  wire [8:0] _T_270 = $signed(_T_269) / 8'sh2; // @[GameLogic.scala 702:66]
  wire [10:0] _GEN_4413 = {{2{_T_270[8]}},_T_270}; // @[GameLogic.scala 702:51]
  wire [10:0] _T_280 = $signed(Ystart_17) + $signed(_GEN_4413); // @[GameLogic.scala 703:51]
  wire  _T_281 = hp <= 4'h0; // @[GameLogic.scala 330:13]
  wire  _T_282 = cngCnt == 4'h0; // @[GameLogic.scala 333:40]
  wire  _T_283 = cngCnt == 4'h1; // @[GameLogic.scala 334:40]
  wire  _T_284 = cngCnt == 4'h2; // @[GameLogic.scala 335:40]
  wire  _GEN_4 = _T_281 & _T_282; // @[GameLogic.scala 330:21]
  wire  _GEN_5 = _T_281 & _T_283; // @[GameLogic.scala 330:21]
  wire  _GEN_6 = _T_281 & _T_284; // @[GameLogic.scala 330:21]
  wire [11:0] _T_286 = {{1{Xstart_17[10]}},Xstart_17}; // @[GameLogic.scala 398:44]
  wire [10:0] _T_288 = _T_286[10:0]; // @[GameLogic.scala 398:44]
  wire [11:0] _T_289 = {{1{Ystart_17[10]}},Ystart_17}; // @[GameLogic.scala 399:44]
  wire [10:0] _T_291 = _T_289[10:0]; // @[GameLogic.scala 399:44]
  wire [10:0] _T_294 = $signed(Xstart_17) + 11'sh20; // @[GameLogic.scala 398:44]
  wire [10:0] _T_300 = $signed(Xstart_17) + 11'sh40; // @[GameLogic.scala 398:44]
  wire [10:0] _T_309 = $signed(Ystart_17) + 11'sh20; // @[GameLogic.scala 399:44]
  wire [10:0] _T_327 = $signed(Ystart_17) + 11'sh40; // @[GameLogic.scala 399:44]
  wire  _T_340 = planetHp < 5'h1; // @[GameLogic.scala 405:19]
  wire  _GEN_8 = _T_340 ? 1'h0 : astInteract_0; // @[GameLogic.scala 405:26]
  wire  _GEN_9 = _T_340 ? 1'h0 : spriteVisibleReg_7; // @[GameLogic.scala 405:26]
  wire  _GEN_10 = _T_340 ? 1'h0 : astInteract_1; // @[GameLogic.scala 405:26]
  wire  _GEN_11 = _T_340 ? 1'h0 : spriteVisibleReg_8; // @[GameLogic.scala 405:26]
  wire  _GEN_12 = _T_340 ? 1'h0 : astInteract_2; // @[GameLogic.scala 405:26]
  wire  _GEN_13 = _T_340 ? 1'h0 : spriteVisibleReg_9; // @[GameLogic.scala 405:26]
  wire  _GEN_14 = _T_340 ? 1'h0 : astInteract_3; // @[GameLogic.scala 405:26]
  wire  _GEN_15 = _T_340 ? 1'h0 : spriteVisibleReg_10; // @[GameLogic.scala 405:26]
  wire  _GEN_16 = _T_340 ? 1'h0 : astInteract_4; // @[GameLogic.scala 405:26]
  wire  _GEN_17 = _T_340 ? 1'h0 : spriteVisibleReg_11; // @[GameLogic.scala 405:26]
  wire  _GEN_18 = _T_340 ? 1'h0 : astInteract_5; // @[GameLogic.scala 405:26]
  wire  _GEN_19 = _T_340 ? 1'h0 : spriteVisibleReg_12; // @[GameLogic.scala 405:26]
  wire  _GEN_20 = _T_340 ? 1'h0 : astInteract_6; // @[GameLogic.scala 405:26]
  wire  _GEN_21 = _T_340 ? 1'h0 : spriteVisibleReg_13; // @[GameLogic.scala 405:26]
  wire  _GEN_22 = _T_340 ? 1'h0 : astInteract_7; // @[GameLogic.scala 405:26]
  wire  _GEN_23 = _T_340 ? 1'h0 : spriteVisibleReg_14; // @[GameLogic.scala 405:26]
  wire  _GEN_24 = _T_340 ? 1'h0 : astInteract_8; // @[GameLogic.scala 405:26]
  wire  _GEN_25 = _T_340 ? 1'h0 : spriteVisibleReg_15; // @[GameLogic.scala 405:26]
  wire  _GEN_26 = _T_340 ? 1'h0 : astInteract_9; // @[GameLogic.scala 405:26]
  wire  _GEN_27 = _T_340 ? 1'h0 : spriteVisibleReg_16; // @[GameLogic.scala 405:26]
  wire  _GEN_28 = _T_340 ? 1'h0 : astInteract_10; // @[GameLogic.scala 405:26]
  wire  _GEN_29 = _T_340 ? 1'h0 : spriteVisibleReg_17; // @[GameLogic.scala 405:26]
  wire  _T_341 = 4'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_342 = 4'h1 == stateReg; // @[Conditional.scala 37:30]
  wire [9:0] _T_345 = viewX + 10'h2; // @[GameLogic.scala 721:22]
  wire [10:0] _T_348 = $signed(Xstart_2) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_351 = $signed(Xstart_3) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_354 = $signed(Xstart_4) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_357 = $signed(Xstart_5) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_360 = $signed(Xstart_6) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_363 = $signed(Xstart_7) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_366 = $signed(Xstart_8) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_369 = $signed(Xstart_9) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_372 = $signed(Xstart_10) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_375 = $signed(Xstart_11) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_378 = $signed(Xstart_12) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_381 = $signed(Xstart_13) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_384 = $signed(Xstart_14) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_387 = $signed(Xstart_15) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_390 = $signed(Xstart_16) - 11'sh2; // @[GameLogic.scala 730:40]
  wire [10:0] _T_393 = $signed(Xstart_17) - 11'sh2; // @[GameLogic.scala 730:40]
  wire  _T_395 = viewX >= 10'h20; // @[GameLogic.scala 734:18]
  wire [9:0] _T_398 = viewX - 10'h20; // @[GameLogic.scala 736:24]
  wire [9:0] _T_401 = _T_398 + 10'h2; // @[GameLogic.scala 736:43]
  wire [6:0] _T_403 = count1 + 7'h1; // @[GameLogic.scala 740:28]
  wire  _T_404 = 4'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_405 = count1 >= 7'h1a; // @[GameLogic.scala 748:19]
  wire  _T_406 = viewX >= 10'h16; // @[GameLogic.scala 753:18]
  wire  _T_407 = count4 == 8'h1; // @[GameLogic.scala 755:21]
  wire  _T_408 = count3 < 7'h9; // @[GameLogic.scala 756:23]
  wire [2:0] _T_410 = level - 3'h1; // @[GameLogic.scala 757:53]
  wire [5:0] _T_411 = _T_410 * 3'h5; // @[GameLogic.scala 757:60]
  wire [5:0] _T_413 = 6'hc + _T_411; // @[GameLogic.scala 757:44]
  wire [7:0] _GEN_4415 = {{1'd0}, count1}; // @[GameLogic.scala 758:48]
  wire [7:0] _T_415 = 8'h8f - _GEN_4415; // @[GameLogic.scala 758:48]
  wire [12:0] _T_416 = count3 * 7'h28; // @[GameLogic.scala 758:66]
  wire [12:0] _GEN_4416 = {{5'd0}, _T_415}; // @[GameLogic.scala 758:57]
  wire [12:0] _T_418 = _GEN_4416 + _T_416; // @[GameLogic.scala 758:57]
  wire [6:0] _T_420 = count3 + 7'h1; // @[GameLogic.scala 761:30]
  wire [5:0] _GEN_37 = _T_408 ? _T_413 : 6'h0; // @[GameLogic.scala 756:30]
  wire [12:0] _GEN_38 = _T_408 ? _T_418 : 13'h0; // @[GameLogic.scala 756:30]
  wire [6:0] _GEN_40 = _T_408 ? _T_420 : 7'h0; // @[GameLogic.scala 756:30]
  wire [5:0] _GEN_42 = _T_407 ? _GEN_37 : 6'h0; // @[GameLogic.scala 755:30]
  wire [12:0] _GEN_43 = _T_407 ? _GEN_38 : 13'h0; // @[GameLogic.scala 755:30]
  wire  _GEN_44 = _T_407 & _T_408; // @[GameLogic.scala 755:30]
  wire [5:0] _GEN_47 = _T_406 ? _GEN_42 : 6'h0; // @[GameLogic.scala 753:27]
  wire [12:0] _GEN_48 = _T_406 ? _GEN_43 : 13'h0; // @[GameLogic.scala 753:27]
  wire  _GEN_49 = _T_406 & _GEN_44; // @[GameLogic.scala 753:27]
  wire  _T_421 = viewX < 10'h16; // @[GameLogic.scala 770:19]
  wire  _T_422 = viewX >= 10'hb; // @[GameLogic.scala 770:37]
  wire  _T_423 = _T_421 & _T_422; // @[GameLogic.scala 770:27]
  wire [5:0] _T_429 = 6'hb + _T_411; // @[GameLogic.scala 773:42]
  wire [5:0] _GEN_52 = _T_408 ? _T_429 : _GEN_47; // @[GameLogic.scala 772:28]
  wire [12:0] _GEN_53 = _T_408 ? _T_418 : _GEN_48; // @[GameLogic.scala 772:28]
  wire  _GEN_54 = _T_408 | _GEN_49; // @[GameLogic.scala 772:28]
  wire [5:0] _GEN_57 = _T_423 ? _GEN_52 : _GEN_47; // @[GameLogic.scala 770:47]
  wire [12:0] _GEN_58 = _T_423 ? _GEN_53 : _GEN_48; // @[GameLogic.scala 770:47]
  wire  _GEN_59 = _T_423 ? _GEN_54 : _GEN_49; // @[GameLogic.scala 770:47]
  wire  _T_437 = viewX < 10'hb; // @[GameLogic.scala 784:18]
  wire [5:0] _T_443 = 6'ha + _T_411; // @[GameLogic.scala 787:42]
  wire [5:0] _GEN_62 = _T_408 ? _T_443 : _GEN_57; // @[GameLogic.scala 786:28]
  wire [12:0] _GEN_63 = _T_408 ? _T_418 : _GEN_58; // @[GameLogic.scala 786:28]
  wire  _GEN_64 = _T_408 | _GEN_59; // @[GameLogic.scala 786:28]
  wire [5:0] _GEN_67 = _T_437 ? _GEN_62 : _GEN_57; // @[GameLogic.scala 784:26]
  wire [12:0] _GEN_68 = _T_437 ? _GEN_63 : _GEN_58; // @[GameLogic.scala 784:26]
  wire  _GEN_69 = _T_437 ? _GEN_64 : _GEN_59; // @[GameLogic.scala 784:26]
  wire  _T_451 = 4'h3 == stateReg; // @[Conditional.scala 37:30]
  wire [5:0] _T_464 = 6'he + _T_411; // @[GameLogic.scala 809:42]
  wire [7:0] _T_466 = 8'h90 - _GEN_4415; // @[GameLogic.scala 810:46]
  wire [12:0] _GEN_4422 = {{5'd0}, _T_466}; // @[GameLogic.scala 810:55]
  wire [12:0] _T_469 = _GEN_4422 + _T_416; // @[GameLogic.scala 810:55]
  wire [5:0] _GEN_76 = _T_408 ? _T_464 : 6'h0; // @[GameLogic.scala 808:28]
  wire [12:0] _GEN_77 = _T_408 ? _T_469 : 13'h0; // @[GameLogic.scala 808:28]
  wire [5:0] _GEN_82 = _T_423 ? _GEN_76 : 6'h0; // @[GameLogic.scala 807:47]
  wire [12:0] _GEN_83 = _T_423 ? _GEN_77 : 13'h0; // @[GameLogic.scala 807:47]
  wire  _GEN_84 = _T_423 & _T_408; // @[GameLogic.scala 807:47]
  wire [5:0] _T_478 = 6'hd + _T_411; // @[GameLogic.scala 822:42]
  wire [5:0] _GEN_88 = _T_408 ? _T_478 : _GEN_82; // @[GameLogic.scala 821:28]
  wire [12:0] _GEN_89 = _T_408 ? _T_469 : _GEN_83; // @[GameLogic.scala 821:28]
  wire  _GEN_90 = _T_408 | _GEN_84; // @[GameLogic.scala 821:28]
  wire [5:0] _GEN_93 = _T_437 ? _GEN_88 : _GEN_82; // @[GameLogic.scala 820:26]
  wire [12:0] _GEN_94 = _T_437 ? _GEN_89 : _GEN_83; // @[GameLogic.scala 820:26]
  wire  _GEN_95 = _T_437 ? _GEN_90 : _GEN_84; // @[GameLogic.scala 820:26]
  wire  _T_486 = 4'h4 == stateReg; // @[Conditional.scala 37:30]
  wire [7:0] _T_494 = 8'h91 - _GEN_4415; // @[GameLogic.scala 837:44]
  wire [12:0] _GEN_4426 = {{5'd0}, _T_494}; // @[GameLogic.scala 837:53]
  wire [12:0] _T_497 = _GEN_4426 + _T_416; // @[GameLogic.scala 837:53]
  wire  _T_500 = planetHp <= 5'h0; // @[GameLogic.scala 841:27]
  wire  _T_501 = level >= 3'h4; // @[GameLogic.scala 845:31]
  wire  _T_502 = $signed(secCnt) >= 8'sha; // @[GameLogic.scala 845:48]
  wire  _T_503 = _T_501 & _T_502; // @[GameLogic.scala 845:38]
  wire [12:0] _GEN_101 = _T_408 ? _T_497 : 13'h0; // @[GameLogic.scala 835:26]
  wire  _T_505 = 4'h5 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_506 = level < 3'h4; // @[GameLogic.scala 850:27]
  wire  _T_507 = start & _T_506; // @[GameLogic.scala 850:18]
  wire [10:0] _T_510 = $signed(Xstart_7) - 11'sh4; // @[GameLogic.scala 294:44]
  wire  _T_511 = planetHp >= 5'h1; // @[GameLogic.scala 295:19]
  wire  _T_512 = $signed(Xstart_7) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_513 = $signed(secCnt) >= 8'sh5; // @[GameLogic.scala 191:45]
  wire  _T_514 = _T_512 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4427 = {{4{Randomizer_1_io_out[6]}},Randomizer_1_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_521 = $signed(_GEN_4427) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire [9:0] _T_522 = viewX; // @[GameLogic.scala 198:47]
  wire [10:0] _GEN_4428 = {{1{_T_522[9]}},_T_522}; // @[GameLogic.scala 198:39]
  wire [10:0] _T_525 = 11'sh2c0 + $signed(_GEN_4428); // @[GameLogic.scala 198:39]
  wire [10:0] _GEN_105 = _T_501 ? $signed(_T_294) : $signed(_T_525); // @[GameLogic.scala 194:26]
  wire  _GEN_107 = _T_514 | _GEN_8; // @[GameLogic.scala 191:53]
  wire  _GEN_108 = _T_514 | _GEN_9; // @[GameLogic.scala 191:53]
  wire  _GEN_115 = kill_0_3 & shotInteract_0; // @[GameLogic.scala 157:41]
  wire  _GEN_116 = kill_0_3 ? shotPop_0 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_117 = kill_0_3 & spriteVisibleReg_2; // @[GameLogic.scala 157:41]
  wire  _GEN_119 = kill_0_0 ? _GEN_115 : shotInteract_0; // @[GameLogic.scala 155:39]
  wire  _GEN_120 = kill_0_0 ? _GEN_116 : shotPop_0; // @[GameLogic.scala 155:39]
  wire  _GEN_121 = kill_0_0 ? _GEN_117 : spriteVisibleReg_2; // @[GameLogic.scala 155:39]
  wire  _GEN_123 = kill_0_3 & shotInteract_1; // @[GameLogic.scala 157:41]
  wire  _GEN_124 = kill_0_3 ? shotPop_1 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_125 = kill_0_3 & spriteVisibleReg_3; // @[GameLogic.scala 157:41]
  wire  _GEN_127 = kill_0_1 ? _GEN_123 : shotInteract_1; // @[GameLogic.scala 155:39]
  wire  _GEN_128 = kill_0_1 ? _GEN_124 : shotPop_1; // @[GameLogic.scala 155:39]
  wire  _GEN_129 = kill_0_1 ? _GEN_125 : spriteVisibleReg_3; // @[GameLogic.scala 155:39]
  wire  _GEN_131 = kill_0_3 & shotInteract_2; // @[GameLogic.scala 157:41]
  wire  _GEN_132 = kill_0_3 ? shotPop_2 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_133 = kill_0_3 & spriteVisibleReg_4; // @[GameLogic.scala 157:41]
  wire  _GEN_135 = kill_0_2 ? _GEN_131 : shotInteract_2; // @[GameLogic.scala 155:39]
  wire  _GEN_136 = kill_0_2 ? _GEN_132 : shotPop_2; // @[GameLogic.scala 155:39]
  wire  _GEN_137 = kill_0_2 ? _GEN_133 : spriteVisibleReg_4; // @[GameLogic.scala 155:39]
  wire  _GEN_139 = kill_0_3 & shotInteract_3; // @[GameLogic.scala 157:41]
  wire  _GEN_140 = kill_0_3 ? shotPop_3 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_141 = kill_0_3 & spriteVisibleReg_5; // @[GameLogic.scala 157:41]
  wire  _GEN_143 = kill_0_3 ? _GEN_139 : shotInteract_3; // @[GameLogic.scala 155:39]
  wire  _GEN_144 = kill_0_3 ? _GEN_140 : shotPop_3; // @[GameLogic.scala 155:39]
  wire  _GEN_145 = kill_0_3 ? _GEN_141 : spriteVisibleReg_5; // @[GameLogic.scala 155:39]
  wire  _GEN_147 = kill_0_3 & shotInteract_4; // @[GameLogic.scala 157:41]
  wire  _GEN_148 = kill_0_3 ? shotPop_4 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_149 = kill_0_3 & spriteVisibleReg_6; // @[GameLogic.scala 157:41]
  wire  _GEN_151 = kill_0_4 ? _GEN_147 : shotInteract_4; // @[GameLogic.scala 155:39]
  wire  _GEN_152 = kill_0_4 ? _GEN_148 : shotPop_4; // @[GameLogic.scala 155:39]
  wire  _GEN_153 = kill_0_4 ? _GEN_149 : spriteVisibleReg_6; // @[GameLogic.scala 155:39]
  wire [10:0] _T_528 = $signed(Xstart_8) - 11'sh4; // @[GameLogic.scala 294:44]
  wire  _T_530 = $signed(Xstart_8) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_532 = _T_530 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4429 = {{4{Randomizer_3_io_out[6]}},Randomizer_3_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_539 = $signed(_GEN_4429) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_157 = _T_532 | _GEN_10; // @[GameLogic.scala 191:53]
  wire  _GEN_158 = _T_532 | _GEN_11; // @[GameLogic.scala 191:53]
  wire  _GEN_165 = kill_1_3 & _GEN_119; // @[GameLogic.scala 157:41]
  wire  _GEN_166 = kill_1_3 ? _GEN_120 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_167 = kill_1_3 & _GEN_121; // @[GameLogic.scala 157:41]
  wire  _GEN_169 = kill_1_0 ? _GEN_165 : _GEN_119; // @[GameLogic.scala 155:39]
  wire  _GEN_170 = kill_1_0 ? _GEN_166 : _GEN_120; // @[GameLogic.scala 155:39]
  wire  _GEN_171 = kill_1_0 ? _GEN_167 : _GEN_121; // @[GameLogic.scala 155:39]
  wire  _GEN_173 = kill_1_3 & _GEN_127; // @[GameLogic.scala 157:41]
  wire  _GEN_174 = kill_1_3 ? _GEN_128 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_175 = kill_1_3 & _GEN_129; // @[GameLogic.scala 157:41]
  wire  _GEN_177 = kill_1_1 ? _GEN_173 : _GEN_127; // @[GameLogic.scala 155:39]
  wire  _GEN_178 = kill_1_1 ? _GEN_174 : _GEN_128; // @[GameLogic.scala 155:39]
  wire  _GEN_179 = kill_1_1 ? _GEN_175 : _GEN_129; // @[GameLogic.scala 155:39]
  wire  _GEN_181 = kill_1_3 & _GEN_135; // @[GameLogic.scala 157:41]
  wire  _GEN_182 = kill_1_3 ? _GEN_136 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_183 = kill_1_3 & _GEN_137; // @[GameLogic.scala 157:41]
  wire  _GEN_185 = kill_1_2 ? _GEN_181 : _GEN_135; // @[GameLogic.scala 155:39]
  wire  _GEN_186 = kill_1_2 ? _GEN_182 : _GEN_136; // @[GameLogic.scala 155:39]
  wire  _GEN_187 = kill_1_2 ? _GEN_183 : _GEN_137; // @[GameLogic.scala 155:39]
  wire  _GEN_189 = kill_1_3 & _GEN_143; // @[GameLogic.scala 157:41]
  wire  _GEN_190 = kill_1_3 ? _GEN_144 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_191 = kill_1_3 & _GEN_145; // @[GameLogic.scala 157:41]
  wire  _GEN_193 = kill_1_3 ? _GEN_189 : _GEN_143; // @[GameLogic.scala 155:39]
  wire  _GEN_194 = kill_1_3 ? _GEN_190 : _GEN_144; // @[GameLogic.scala 155:39]
  wire  _GEN_195 = kill_1_3 ? _GEN_191 : _GEN_145; // @[GameLogic.scala 155:39]
  wire  _GEN_197 = kill_1_3 & _GEN_151; // @[GameLogic.scala 157:41]
  wire  _GEN_198 = kill_1_3 ? _GEN_152 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_199 = kill_1_3 & _GEN_153; // @[GameLogic.scala 157:41]
  wire  _GEN_201 = kill_1_4 ? _GEN_197 : _GEN_151; // @[GameLogic.scala 155:39]
  wire  _GEN_202 = kill_1_4 ? _GEN_198 : _GEN_152; // @[GameLogic.scala 155:39]
  wire  _GEN_203 = kill_1_4 ? _GEN_199 : _GEN_153; // @[GameLogic.scala 155:39]
  wire [10:0] _T_546 = $signed(Xstart_9) - 11'sh4; // @[GameLogic.scala 294:44]
  wire  _T_548 = $signed(Xstart_9) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_550 = _T_548 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4431 = {{4{Randomizer_5_io_out[6]}},Randomizer_5_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_557 = $signed(_GEN_4431) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_207 = _T_550 | _GEN_12; // @[GameLogic.scala 191:53]
  wire  _GEN_208 = _T_550 | _GEN_13; // @[GameLogic.scala 191:53]
  wire  _GEN_215 = kill_2_3 & _GEN_169; // @[GameLogic.scala 157:41]
  wire  _GEN_216 = kill_2_3 ? _GEN_170 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_217 = kill_2_3 & _GEN_171; // @[GameLogic.scala 157:41]
  wire  _GEN_219 = kill_2_0 ? _GEN_215 : _GEN_169; // @[GameLogic.scala 155:39]
  wire  _GEN_220 = kill_2_0 ? _GEN_216 : _GEN_170; // @[GameLogic.scala 155:39]
  wire  _GEN_221 = kill_2_0 ? _GEN_217 : _GEN_171; // @[GameLogic.scala 155:39]
  wire  _GEN_223 = kill_2_3 & _GEN_177; // @[GameLogic.scala 157:41]
  wire  _GEN_224 = kill_2_3 ? _GEN_178 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_225 = kill_2_3 & _GEN_179; // @[GameLogic.scala 157:41]
  wire  _GEN_227 = kill_2_1 ? _GEN_223 : _GEN_177; // @[GameLogic.scala 155:39]
  wire  _GEN_228 = kill_2_1 ? _GEN_224 : _GEN_178; // @[GameLogic.scala 155:39]
  wire  _GEN_229 = kill_2_1 ? _GEN_225 : _GEN_179; // @[GameLogic.scala 155:39]
  wire  _GEN_231 = kill_2_3 & _GEN_185; // @[GameLogic.scala 157:41]
  wire  _GEN_232 = kill_2_3 ? _GEN_186 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_233 = kill_2_3 & _GEN_187; // @[GameLogic.scala 157:41]
  wire  _GEN_235 = kill_2_2 ? _GEN_231 : _GEN_185; // @[GameLogic.scala 155:39]
  wire  _GEN_236 = kill_2_2 ? _GEN_232 : _GEN_186; // @[GameLogic.scala 155:39]
  wire  _GEN_237 = kill_2_2 ? _GEN_233 : _GEN_187; // @[GameLogic.scala 155:39]
  wire  _GEN_239 = kill_2_3 & _GEN_193; // @[GameLogic.scala 157:41]
  wire  _GEN_240 = kill_2_3 ? _GEN_194 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_241 = kill_2_3 & _GEN_195; // @[GameLogic.scala 157:41]
  wire  _GEN_243 = kill_2_3 ? _GEN_239 : _GEN_193; // @[GameLogic.scala 155:39]
  wire  _GEN_244 = kill_2_3 ? _GEN_240 : _GEN_194; // @[GameLogic.scala 155:39]
  wire  _GEN_245 = kill_2_3 ? _GEN_241 : _GEN_195; // @[GameLogic.scala 155:39]
  wire  _GEN_247 = kill_2_3 & _GEN_201; // @[GameLogic.scala 157:41]
  wire  _GEN_248 = kill_2_3 ? _GEN_202 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_249 = kill_2_3 & _GEN_203; // @[GameLogic.scala 157:41]
  wire  _GEN_251 = kill_2_4 ? _GEN_247 : _GEN_201; // @[GameLogic.scala 155:39]
  wire  _GEN_252 = kill_2_4 ? _GEN_248 : _GEN_202; // @[GameLogic.scala 155:39]
  wire  _GEN_253 = kill_2_4 ? _GEN_249 : _GEN_203; // @[GameLogic.scala 155:39]
  wire  _T_562 = level >= 3'h1; // @[GameLogic.scala 854:31]
  wire  _T_565 = _T_501 & _T_513; // @[GameLogic.scala 854:56]
  wire  _GEN_259 = _T_507 ? _GEN_219 : shotInteract_0; // @[GameLogic.scala 850:34]
  wire  _GEN_260 = _T_507 ? _GEN_220 : shotPop_0; // @[GameLogic.scala 850:34]
  wire  _GEN_261 = _T_507 ? _GEN_221 : spriteVisibleReg_2; // @[GameLogic.scala 850:34]
  wire  _GEN_262 = _T_507 ? _GEN_227 : shotInteract_1; // @[GameLogic.scala 850:34]
  wire  _GEN_263 = _T_507 ? _GEN_228 : shotPop_1; // @[GameLogic.scala 850:34]
  wire  _GEN_264 = _T_507 ? _GEN_229 : spriteVisibleReg_3; // @[GameLogic.scala 850:34]
  wire  _GEN_265 = _T_507 ? _GEN_235 : shotInteract_2; // @[GameLogic.scala 850:34]
  wire  _GEN_266 = _T_507 ? _GEN_236 : shotPop_2; // @[GameLogic.scala 850:34]
  wire  _GEN_267 = _T_507 ? _GEN_237 : spriteVisibleReg_4; // @[GameLogic.scala 850:34]
  wire  _GEN_268 = _T_507 ? _GEN_243 : shotInteract_3; // @[GameLogic.scala 850:34]
  wire  _GEN_269 = _T_507 ? _GEN_244 : shotPop_3; // @[GameLogic.scala 850:34]
  wire  _GEN_270 = _T_507 ? _GEN_245 : spriteVisibleReg_5; // @[GameLogic.scala 850:34]
  wire  _GEN_271 = _T_507 ? _GEN_251 : shotInteract_4; // @[GameLogic.scala 850:34]
  wire  _GEN_272 = _T_507 ? _GEN_252 : shotPop_4; // @[GameLogic.scala 850:34]
  wire  _GEN_273 = _T_507 ? _GEN_253 : spriteVisibleReg_6; // @[GameLogic.scala 850:34]
  wire  _T_570 = 4'h6 == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_573 = $signed(Xstart_10) - 11'sh4; // @[GameLogic.scala 294:44]
  wire  _T_575 = $signed(Xstart_10) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_577 = _T_575 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4433 = {{4{Randomizer_7_io_out[6]}},Randomizer_7_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_584 = $signed(_GEN_4433) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_285 = _T_577 | _GEN_14; // @[GameLogic.scala 191:53]
  wire  _GEN_286 = _T_577 | _GEN_15; // @[GameLogic.scala 191:53]
  wire  _GEN_293 = kill_3_3 & shotInteract_0; // @[GameLogic.scala 157:41]
  wire  _GEN_294 = kill_3_3 ? shotPop_0 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_295 = kill_3_3 & spriteVisibleReg_2; // @[GameLogic.scala 157:41]
  wire  _GEN_297 = kill_3_0 ? _GEN_293 : shotInteract_0; // @[GameLogic.scala 155:39]
  wire  _GEN_298 = kill_3_0 ? _GEN_294 : shotPop_0; // @[GameLogic.scala 155:39]
  wire  _GEN_299 = kill_3_0 ? _GEN_295 : spriteVisibleReg_2; // @[GameLogic.scala 155:39]
  wire  _GEN_301 = kill_3_3 & shotInteract_1; // @[GameLogic.scala 157:41]
  wire  _GEN_302 = kill_3_3 ? shotPop_1 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_303 = kill_3_3 & spriteVisibleReg_3; // @[GameLogic.scala 157:41]
  wire  _GEN_305 = kill_3_1 ? _GEN_301 : shotInteract_1; // @[GameLogic.scala 155:39]
  wire  _GEN_306 = kill_3_1 ? _GEN_302 : shotPop_1; // @[GameLogic.scala 155:39]
  wire  _GEN_307 = kill_3_1 ? _GEN_303 : spriteVisibleReg_3; // @[GameLogic.scala 155:39]
  wire  _GEN_309 = kill_3_3 & shotInteract_2; // @[GameLogic.scala 157:41]
  wire  _GEN_310 = kill_3_3 ? shotPop_2 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_311 = kill_3_3 & spriteVisibleReg_4; // @[GameLogic.scala 157:41]
  wire  _GEN_313 = kill_3_2 ? _GEN_309 : shotInteract_2; // @[GameLogic.scala 155:39]
  wire  _GEN_314 = kill_3_2 ? _GEN_310 : shotPop_2; // @[GameLogic.scala 155:39]
  wire  _GEN_315 = kill_3_2 ? _GEN_311 : spriteVisibleReg_4; // @[GameLogic.scala 155:39]
  wire  _GEN_317 = kill_3_3 & shotInteract_3; // @[GameLogic.scala 157:41]
  wire  _GEN_318 = kill_3_3 ? shotPop_3 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_319 = kill_3_3 & spriteVisibleReg_5; // @[GameLogic.scala 157:41]
  wire  _GEN_321 = kill_3_3 ? _GEN_317 : shotInteract_3; // @[GameLogic.scala 155:39]
  wire  _GEN_322 = kill_3_3 ? _GEN_318 : shotPop_3; // @[GameLogic.scala 155:39]
  wire  _GEN_323 = kill_3_3 ? _GEN_319 : spriteVisibleReg_5; // @[GameLogic.scala 155:39]
  wire  _GEN_325 = kill_3_3 & shotInteract_4; // @[GameLogic.scala 157:41]
  wire  _GEN_326 = kill_3_3 ? shotPop_4 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_327 = kill_3_3 & spriteVisibleReg_6; // @[GameLogic.scala 157:41]
  wire  _GEN_329 = kill_3_4 ? _GEN_325 : shotInteract_4; // @[GameLogic.scala 155:39]
  wire  _GEN_330 = kill_3_4 ? _GEN_326 : shotPop_4; // @[GameLogic.scala 155:39]
  wire  _GEN_331 = kill_3_4 ? _GEN_327 : spriteVisibleReg_6; // @[GameLogic.scala 155:39]
  wire [10:0] _T_591 = $signed(Xstart_11) - 11'sh5; // @[GameLogic.scala 294:44]
  wire  _T_593 = $signed(Xstart_11) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_595 = _T_593 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4435 = {{4{Randomizer_9_io_out[6]}},Randomizer_9_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_602 = $signed(_GEN_4435) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_335 = _T_595 | _GEN_16; // @[GameLogic.scala 191:53]
  wire  _GEN_336 = _T_595 | _GEN_17; // @[GameLogic.scala 191:53]
  wire  _GEN_343 = kill_4_3 & _GEN_297; // @[GameLogic.scala 157:41]
  wire  _GEN_344 = kill_4_3 ? _GEN_298 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_345 = kill_4_3 & _GEN_299; // @[GameLogic.scala 157:41]
  wire  _GEN_347 = kill_4_0 ? _GEN_343 : _GEN_297; // @[GameLogic.scala 155:39]
  wire  _GEN_348 = kill_4_0 ? _GEN_344 : _GEN_298; // @[GameLogic.scala 155:39]
  wire  _GEN_349 = kill_4_0 ? _GEN_345 : _GEN_299; // @[GameLogic.scala 155:39]
  wire  _GEN_351 = kill_4_3 & _GEN_305; // @[GameLogic.scala 157:41]
  wire  _GEN_352 = kill_4_3 ? _GEN_306 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_353 = kill_4_3 & _GEN_307; // @[GameLogic.scala 157:41]
  wire  _GEN_355 = kill_4_1 ? _GEN_351 : _GEN_305; // @[GameLogic.scala 155:39]
  wire  _GEN_356 = kill_4_1 ? _GEN_352 : _GEN_306; // @[GameLogic.scala 155:39]
  wire  _GEN_357 = kill_4_1 ? _GEN_353 : _GEN_307; // @[GameLogic.scala 155:39]
  wire  _GEN_359 = kill_4_3 & _GEN_313; // @[GameLogic.scala 157:41]
  wire  _GEN_360 = kill_4_3 ? _GEN_314 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_361 = kill_4_3 & _GEN_315; // @[GameLogic.scala 157:41]
  wire  _GEN_363 = kill_4_2 ? _GEN_359 : _GEN_313; // @[GameLogic.scala 155:39]
  wire  _GEN_364 = kill_4_2 ? _GEN_360 : _GEN_314; // @[GameLogic.scala 155:39]
  wire  _GEN_365 = kill_4_2 ? _GEN_361 : _GEN_315; // @[GameLogic.scala 155:39]
  wire  _GEN_367 = kill_4_3 & _GEN_321; // @[GameLogic.scala 157:41]
  wire  _GEN_368 = kill_4_3 ? _GEN_322 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_369 = kill_4_3 & _GEN_323; // @[GameLogic.scala 157:41]
  wire  _GEN_371 = kill_4_3 ? _GEN_367 : _GEN_321; // @[GameLogic.scala 155:39]
  wire  _GEN_372 = kill_4_3 ? _GEN_368 : _GEN_322; // @[GameLogic.scala 155:39]
  wire  _GEN_373 = kill_4_3 ? _GEN_369 : _GEN_323; // @[GameLogic.scala 155:39]
  wire  _GEN_375 = kill_4_3 & _GEN_329; // @[GameLogic.scala 157:41]
  wire  _GEN_376 = kill_4_3 ? _GEN_330 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_377 = kill_4_3 & _GEN_331; // @[GameLogic.scala 157:41]
  wire  _GEN_379 = kill_4_4 ? _GEN_375 : _GEN_329; // @[GameLogic.scala 155:39]
  wire  _GEN_380 = kill_4_4 ? _GEN_376 : _GEN_330; // @[GameLogic.scala 155:39]
  wire  _GEN_381 = kill_4_4 ? _GEN_377 : _GEN_331; // @[GameLogic.scala 155:39]
  wire [10:0] _T_609 = $signed(Xstart_12) - 11'sh5; // @[GameLogic.scala 294:44]
  wire  _T_611 = $signed(Xstart_12) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_613 = _T_611 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4437 = {{4{Randomizer_11_io_out[6]}},Randomizer_11_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_620 = $signed(_GEN_4437) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_385 = _T_613 | _GEN_18; // @[GameLogic.scala 191:53]
  wire  _GEN_386 = _T_613 | _GEN_19; // @[GameLogic.scala 191:53]
  wire  _GEN_393 = kill_5_3 & _GEN_347; // @[GameLogic.scala 157:41]
  wire  _GEN_394 = kill_5_3 ? _GEN_348 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_395 = kill_5_3 & _GEN_349; // @[GameLogic.scala 157:41]
  wire  _GEN_397 = kill_5_0 ? _GEN_393 : _GEN_347; // @[GameLogic.scala 155:39]
  wire  _GEN_398 = kill_5_0 ? _GEN_394 : _GEN_348; // @[GameLogic.scala 155:39]
  wire  _GEN_399 = kill_5_0 ? _GEN_395 : _GEN_349; // @[GameLogic.scala 155:39]
  wire  _GEN_401 = kill_5_3 & _GEN_355; // @[GameLogic.scala 157:41]
  wire  _GEN_402 = kill_5_3 ? _GEN_356 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_403 = kill_5_3 & _GEN_357; // @[GameLogic.scala 157:41]
  wire  _GEN_405 = kill_5_1 ? _GEN_401 : _GEN_355; // @[GameLogic.scala 155:39]
  wire  _GEN_406 = kill_5_1 ? _GEN_402 : _GEN_356; // @[GameLogic.scala 155:39]
  wire  _GEN_407 = kill_5_1 ? _GEN_403 : _GEN_357; // @[GameLogic.scala 155:39]
  wire  _GEN_409 = kill_5_3 & _GEN_363; // @[GameLogic.scala 157:41]
  wire  _GEN_410 = kill_5_3 ? _GEN_364 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_411 = kill_5_3 & _GEN_365; // @[GameLogic.scala 157:41]
  wire  _GEN_413 = kill_5_2 ? _GEN_409 : _GEN_363; // @[GameLogic.scala 155:39]
  wire  _GEN_414 = kill_5_2 ? _GEN_410 : _GEN_364; // @[GameLogic.scala 155:39]
  wire  _GEN_415 = kill_5_2 ? _GEN_411 : _GEN_365; // @[GameLogic.scala 155:39]
  wire  _GEN_417 = kill_5_3 & _GEN_371; // @[GameLogic.scala 157:41]
  wire  _GEN_418 = kill_5_3 ? _GEN_372 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_419 = kill_5_3 & _GEN_373; // @[GameLogic.scala 157:41]
  wire  _GEN_421 = kill_5_3 ? _GEN_417 : _GEN_371; // @[GameLogic.scala 155:39]
  wire  _GEN_422 = kill_5_3 ? _GEN_418 : _GEN_372; // @[GameLogic.scala 155:39]
  wire  _GEN_423 = kill_5_3 ? _GEN_419 : _GEN_373; // @[GameLogic.scala 155:39]
  wire  _GEN_425 = kill_5_3 & _GEN_379; // @[GameLogic.scala 157:41]
  wire  _GEN_426 = kill_5_3 ? _GEN_380 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_427 = kill_5_3 & _GEN_381; // @[GameLogic.scala 157:41]
  wire  _GEN_429 = kill_5_4 ? _GEN_425 : _GEN_379; // @[GameLogic.scala 155:39]
  wire  _GEN_430 = kill_5_4 ? _GEN_426 : _GEN_380; // @[GameLogic.scala 155:39]
  wire  _GEN_431 = kill_5_4 ? _GEN_427 : _GEN_381; // @[GameLogic.scala 155:39]
  wire  _T_625 = level >= 3'h2; // @[GameLogic.scala 865:29]
  wire  _T_627 = 4'h7 == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_630 = $signed(Xstart_13) - 11'sh5; // @[GameLogic.scala 294:44]
  wire  _T_632 = $signed(Xstart_13) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_634 = _T_632 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4439 = {{4{Randomizer_13_io_out[6]}},Randomizer_13_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_641 = $signed(_GEN_4439) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_435 = _T_634 | _GEN_20; // @[GameLogic.scala 191:53]
  wire  _GEN_436 = _T_634 | _GEN_21; // @[GameLogic.scala 191:53]
  wire  _GEN_443 = kill_6_3 & shotInteract_0; // @[GameLogic.scala 157:41]
  wire  _GEN_444 = kill_6_3 ? shotPop_0 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_445 = kill_6_3 & spriteVisibleReg_2; // @[GameLogic.scala 157:41]
  wire  _GEN_447 = kill_6_0 ? _GEN_443 : shotInteract_0; // @[GameLogic.scala 155:39]
  wire  _GEN_448 = kill_6_0 ? _GEN_444 : shotPop_0; // @[GameLogic.scala 155:39]
  wire  _GEN_449 = kill_6_0 ? _GEN_445 : spriteVisibleReg_2; // @[GameLogic.scala 155:39]
  wire  _GEN_451 = kill_6_3 & shotInteract_1; // @[GameLogic.scala 157:41]
  wire  _GEN_452 = kill_6_3 ? shotPop_1 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_453 = kill_6_3 & spriteVisibleReg_3; // @[GameLogic.scala 157:41]
  wire  _GEN_455 = kill_6_1 ? _GEN_451 : shotInteract_1; // @[GameLogic.scala 155:39]
  wire  _GEN_456 = kill_6_1 ? _GEN_452 : shotPop_1; // @[GameLogic.scala 155:39]
  wire  _GEN_457 = kill_6_1 ? _GEN_453 : spriteVisibleReg_3; // @[GameLogic.scala 155:39]
  wire  _GEN_459 = kill_6_3 & shotInteract_2; // @[GameLogic.scala 157:41]
  wire  _GEN_460 = kill_6_3 ? shotPop_2 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_461 = kill_6_3 & spriteVisibleReg_4; // @[GameLogic.scala 157:41]
  wire  _GEN_463 = kill_6_2 ? _GEN_459 : shotInteract_2; // @[GameLogic.scala 155:39]
  wire  _GEN_464 = kill_6_2 ? _GEN_460 : shotPop_2; // @[GameLogic.scala 155:39]
  wire  _GEN_465 = kill_6_2 ? _GEN_461 : spriteVisibleReg_4; // @[GameLogic.scala 155:39]
  wire  _GEN_467 = kill_6_3 & shotInteract_3; // @[GameLogic.scala 157:41]
  wire  _GEN_468 = kill_6_3 ? shotPop_3 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_469 = kill_6_3 & spriteVisibleReg_5; // @[GameLogic.scala 157:41]
  wire  _GEN_471 = kill_6_3 ? _GEN_467 : shotInteract_3; // @[GameLogic.scala 155:39]
  wire  _GEN_472 = kill_6_3 ? _GEN_468 : shotPop_3; // @[GameLogic.scala 155:39]
  wire  _GEN_473 = kill_6_3 ? _GEN_469 : spriteVisibleReg_5; // @[GameLogic.scala 155:39]
  wire  _GEN_475 = kill_6_3 & shotInteract_4; // @[GameLogic.scala 157:41]
  wire  _GEN_476 = kill_6_3 ? shotPop_4 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_477 = kill_6_3 & spriteVisibleReg_6; // @[GameLogic.scala 157:41]
  wire  _GEN_479 = kill_6_4 ? _GEN_475 : shotInteract_4; // @[GameLogic.scala 155:39]
  wire  _GEN_480 = kill_6_4 ? _GEN_476 : shotPop_4; // @[GameLogic.scala 155:39]
  wire  _GEN_481 = kill_6_4 ? _GEN_477 : spriteVisibleReg_6; // @[GameLogic.scala 155:39]
  wire [10:0] _T_648 = $signed(Xstart_14) - 11'sh3; // @[GameLogic.scala 294:44]
  wire  _T_650 = $signed(Xstart_14) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_652 = _T_650 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4441 = {{4{Randomizer_15_io_out[6]}},Randomizer_15_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_659 = $signed(_GEN_4441) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_485 = _T_652 | _GEN_22; // @[GameLogic.scala 191:53]
  wire  _GEN_486 = _T_652 | _GEN_23; // @[GameLogic.scala 191:53]
  wire  _GEN_493 = kill_7_3 & _GEN_447; // @[GameLogic.scala 157:41]
  wire  _GEN_494 = kill_7_3 ? _GEN_448 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_495 = kill_7_3 & _GEN_449; // @[GameLogic.scala 157:41]
  wire  _GEN_497 = kill_7_0 ? _GEN_493 : _GEN_447; // @[GameLogic.scala 155:39]
  wire  _GEN_498 = kill_7_0 ? _GEN_494 : _GEN_448; // @[GameLogic.scala 155:39]
  wire  _GEN_499 = kill_7_0 ? _GEN_495 : _GEN_449; // @[GameLogic.scala 155:39]
  wire  _GEN_501 = kill_7_3 & _GEN_455; // @[GameLogic.scala 157:41]
  wire  _GEN_502 = kill_7_3 ? _GEN_456 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_503 = kill_7_3 & _GEN_457; // @[GameLogic.scala 157:41]
  wire  _GEN_505 = kill_7_1 ? _GEN_501 : _GEN_455; // @[GameLogic.scala 155:39]
  wire  _GEN_506 = kill_7_1 ? _GEN_502 : _GEN_456; // @[GameLogic.scala 155:39]
  wire  _GEN_507 = kill_7_1 ? _GEN_503 : _GEN_457; // @[GameLogic.scala 155:39]
  wire  _GEN_509 = kill_7_3 & _GEN_463; // @[GameLogic.scala 157:41]
  wire  _GEN_510 = kill_7_3 ? _GEN_464 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_511 = kill_7_3 & _GEN_465; // @[GameLogic.scala 157:41]
  wire  _GEN_513 = kill_7_2 ? _GEN_509 : _GEN_463; // @[GameLogic.scala 155:39]
  wire  _GEN_514 = kill_7_2 ? _GEN_510 : _GEN_464; // @[GameLogic.scala 155:39]
  wire  _GEN_515 = kill_7_2 ? _GEN_511 : _GEN_465; // @[GameLogic.scala 155:39]
  wire  _GEN_517 = kill_7_3 & _GEN_471; // @[GameLogic.scala 157:41]
  wire  _GEN_518 = kill_7_3 ? _GEN_472 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_519 = kill_7_3 & _GEN_473; // @[GameLogic.scala 157:41]
  wire  _GEN_521 = kill_7_3 ? _GEN_517 : _GEN_471; // @[GameLogic.scala 155:39]
  wire  _GEN_522 = kill_7_3 ? _GEN_518 : _GEN_472; // @[GameLogic.scala 155:39]
  wire  _GEN_523 = kill_7_3 ? _GEN_519 : _GEN_473; // @[GameLogic.scala 155:39]
  wire  _GEN_525 = kill_7_3 & _GEN_479; // @[GameLogic.scala 157:41]
  wire  _GEN_526 = kill_7_3 ? _GEN_480 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_527 = kill_7_3 & _GEN_481; // @[GameLogic.scala 157:41]
  wire  _GEN_529 = kill_7_4 ? _GEN_525 : _GEN_479; // @[GameLogic.scala 155:39]
  wire  _GEN_530 = kill_7_4 ? _GEN_526 : _GEN_480; // @[GameLogic.scala 155:39]
  wire  _GEN_531 = kill_7_4 ? _GEN_527 : _GEN_481; // @[GameLogic.scala 155:39]
  wire [10:0] _T_666 = $signed(Xstart_15) - 11'sh3; // @[GameLogic.scala 294:44]
  wire  _T_668 = $signed(Xstart_15) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_670 = _T_668 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4443 = {{4{Randomizer_17_io_out[6]}},Randomizer_17_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_677 = $signed(_GEN_4443) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_535 = _T_670 | _GEN_24; // @[GameLogic.scala 191:53]
  wire  _GEN_536 = _T_670 | _GEN_25; // @[GameLogic.scala 191:53]
  wire  _GEN_543 = kill_8_3 & _GEN_497; // @[GameLogic.scala 157:41]
  wire  _GEN_544 = kill_8_3 ? _GEN_498 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_545 = kill_8_3 & _GEN_499; // @[GameLogic.scala 157:41]
  wire  _GEN_547 = kill_8_0 ? _GEN_543 : _GEN_497; // @[GameLogic.scala 155:39]
  wire  _GEN_548 = kill_8_0 ? _GEN_544 : _GEN_498; // @[GameLogic.scala 155:39]
  wire  _GEN_549 = kill_8_0 ? _GEN_545 : _GEN_499; // @[GameLogic.scala 155:39]
  wire  _GEN_551 = kill_8_3 & _GEN_505; // @[GameLogic.scala 157:41]
  wire  _GEN_552 = kill_8_3 ? _GEN_506 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_553 = kill_8_3 & _GEN_507; // @[GameLogic.scala 157:41]
  wire  _GEN_555 = kill_8_1 ? _GEN_551 : _GEN_505; // @[GameLogic.scala 155:39]
  wire  _GEN_556 = kill_8_1 ? _GEN_552 : _GEN_506; // @[GameLogic.scala 155:39]
  wire  _GEN_557 = kill_8_1 ? _GEN_553 : _GEN_507; // @[GameLogic.scala 155:39]
  wire  _GEN_559 = kill_8_3 & _GEN_513; // @[GameLogic.scala 157:41]
  wire  _GEN_560 = kill_8_3 ? _GEN_514 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_561 = kill_8_3 & _GEN_515; // @[GameLogic.scala 157:41]
  wire  _GEN_563 = kill_8_2 ? _GEN_559 : _GEN_513; // @[GameLogic.scala 155:39]
  wire  _GEN_564 = kill_8_2 ? _GEN_560 : _GEN_514; // @[GameLogic.scala 155:39]
  wire  _GEN_565 = kill_8_2 ? _GEN_561 : _GEN_515; // @[GameLogic.scala 155:39]
  wire  _GEN_567 = kill_8_3 & _GEN_521; // @[GameLogic.scala 157:41]
  wire  _GEN_568 = kill_8_3 ? _GEN_522 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_569 = kill_8_3 & _GEN_523; // @[GameLogic.scala 157:41]
  wire  _GEN_571 = kill_8_3 ? _GEN_567 : _GEN_521; // @[GameLogic.scala 155:39]
  wire  _GEN_572 = kill_8_3 ? _GEN_568 : _GEN_522; // @[GameLogic.scala 155:39]
  wire  _GEN_573 = kill_8_3 ? _GEN_569 : _GEN_523; // @[GameLogic.scala 155:39]
  wire  _GEN_575 = kill_8_3 & _GEN_529; // @[GameLogic.scala 157:41]
  wire  _GEN_576 = kill_8_3 ? _GEN_530 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_577 = kill_8_3 & _GEN_531; // @[GameLogic.scala 157:41]
  wire  _GEN_579 = kill_8_4 ? _GEN_575 : _GEN_529; // @[GameLogic.scala 155:39]
  wire  _GEN_580 = kill_8_4 ? _GEN_576 : _GEN_530; // @[GameLogic.scala 155:39]
  wire  _GEN_581 = kill_8_4 ? _GEN_577 : _GEN_531; // @[GameLogic.scala 155:39]
  wire  _T_682 = level >= 3'h3; // @[GameLogic.scala 872:29]
  wire  _T_684 = 4'h8 == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_687 = $signed(Xstart_16) - 11'sh4; // @[GameLogic.scala 169:44]
  wire  _T_688 = planetHp > 5'h0; // @[GameLogic.scala 170:19]
  wire  _T_689 = $signed(Xstart_16) <= 11'sh2; // @[GameLogic.scala 191:28]
  wire  _T_691 = _T_689 & _T_513; // @[GameLogic.scala 191:35]
  wire [10:0] _GEN_4445 = {{4{Randomizer_19_io_out[6]}},Randomizer_19_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_698 = $signed(_GEN_4445) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_585 = _T_691 | _GEN_26; // @[GameLogic.scala 191:53]
  wire  _GEN_586 = _T_691 | _GEN_27; // @[GameLogic.scala 191:53]
  wire  _GEN_593 = kill_9_0 ? 1'h0 : shotInteract_0; // @[GameLogic.scala 174:39]
  wire  _GEN_594 = kill_9_0 | shotPop_0; // @[GameLogic.scala 174:39]
  wire  _GEN_595 = kill_9_0 ? 1'h0 : spriteVisibleReg_2; // @[GameLogic.scala 174:39]
  wire  _GEN_596 = kill_9_1 ? 1'h0 : shotInteract_1; // @[GameLogic.scala 174:39]
  wire  _GEN_597 = kill_9_1 | shotPop_1; // @[GameLogic.scala 174:39]
  wire  _GEN_598 = kill_9_1 ? 1'h0 : spriteVisibleReg_3; // @[GameLogic.scala 174:39]
  wire  _GEN_599 = kill_9_2 ? 1'h0 : shotInteract_2; // @[GameLogic.scala 174:39]
  wire  _GEN_600 = kill_9_2 | shotPop_2; // @[GameLogic.scala 174:39]
  wire  _GEN_601 = kill_9_2 ? 1'h0 : spriteVisibleReg_4; // @[GameLogic.scala 174:39]
  wire  _T_705 = 4'h9 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_706 = $signed(secCnt) >= 8'shb; // @[GameLogic.scala 881:19]
  wire [10:0] _GEN_4447 = {{4{Randomizer_21_io_out[6]}},Randomizer_21_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_720 = $signed(_GEN_4447) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire [10:0] _GEN_4449 = {{4{Randomizer_23_io_out[6]}},Randomizer_23_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_738 = $signed(_GEN_4449) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire [10:0] _GEN_4451 = {{4{Randomizer_25_io_out[6]}},Randomizer_25_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_756 = $signed(_GEN_4451) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire [10:0] _GEN_4453 = {{4{Randomizer_27_io_out[6]}},Randomizer_27_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_774 = $signed(_GEN_4453) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_674 = kill_4_3 & _GEN_219; // @[GameLogic.scala 157:41]
  wire  _GEN_675 = kill_4_3 ? _GEN_220 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_676 = kill_4_3 & _GEN_221; // @[GameLogic.scala 157:41]
  wire  _GEN_678 = kill_4_0 ? _GEN_674 : _GEN_219; // @[GameLogic.scala 155:39]
  wire  _GEN_679 = kill_4_0 ? _GEN_675 : _GEN_220; // @[GameLogic.scala 155:39]
  wire  _GEN_680 = kill_4_0 ? _GEN_676 : _GEN_221; // @[GameLogic.scala 155:39]
  wire  _GEN_682 = kill_4_3 & _GEN_227; // @[GameLogic.scala 157:41]
  wire  _GEN_683 = kill_4_3 ? _GEN_228 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_684 = kill_4_3 & _GEN_229; // @[GameLogic.scala 157:41]
  wire  _GEN_686 = kill_4_1 ? _GEN_682 : _GEN_227; // @[GameLogic.scala 155:39]
  wire  _GEN_687 = kill_4_1 ? _GEN_683 : _GEN_228; // @[GameLogic.scala 155:39]
  wire  _GEN_688 = kill_4_1 ? _GEN_684 : _GEN_229; // @[GameLogic.scala 155:39]
  wire  _GEN_690 = kill_4_3 & _GEN_235; // @[GameLogic.scala 157:41]
  wire  _GEN_691 = kill_4_3 ? _GEN_236 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_692 = kill_4_3 & _GEN_237; // @[GameLogic.scala 157:41]
  wire  _GEN_694 = kill_4_2 ? _GEN_690 : _GEN_235; // @[GameLogic.scala 155:39]
  wire  _GEN_695 = kill_4_2 ? _GEN_691 : _GEN_236; // @[GameLogic.scala 155:39]
  wire  _GEN_696 = kill_4_2 ? _GEN_692 : _GEN_237; // @[GameLogic.scala 155:39]
  wire  _GEN_698 = kill_4_3 & _GEN_243; // @[GameLogic.scala 157:41]
  wire  _GEN_699 = kill_4_3 ? _GEN_244 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_700 = kill_4_3 & _GEN_245; // @[GameLogic.scala 157:41]
  wire  _GEN_702 = kill_4_3 ? _GEN_698 : _GEN_243; // @[GameLogic.scala 155:39]
  wire  _GEN_703 = kill_4_3 ? _GEN_699 : _GEN_244; // @[GameLogic.scala 155:39]
  wire  _GEN_704 = kill_4_3 ? _GEN_700 : _GEN_245; // @[GameLogic.scala 155:39]
  wire  _GEN_706 = kill_4_3 & _GEN_251; // @[GameLogic.scala 157:41]
  wire  _GEN_707 = kill_4_3 ? _GEN_252 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_708 = kill_4_3 & _GEN_253; // @[GameLogic.scala 157:41]
  wire  _GEN_710 = kill_4_4 ? _GEN_706 : _GEN_251; // @[GameLogic.scala 155:39]
  wire  _GEN_711 = kill_4_4 ? _GEN_707 : _GEN_252; // @[GameLogic.scala 155:39]
  wire  _GEN_712 = kill_4_4 ? _GEN_708 : _GEN_253; // @[GameLogic.scala 155:39]
  wire [10:0] _GEN_4455 = {{4{Randomizer_29_io_out[6]}},Randomizer_29_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_792 = $signed(_GEN_4455) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_724 = kill_5_3 & _GEN_678; // @[GameLogic.scala 157:41]
  wire  _GEN_725 = kill_5_3 ? _GEN_679 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_726 = kill_5_3 & _GEN_680; // @[GameLogic.scala 157:41]
  wire  _GEN_728 = kill_5_0 ? _GEN_724 : _GEN_678; // @[GameLogic.scala 155:39]
  wire  _GEN_729 = kill_5_0 ? _GEN_725 : _GEN_679; // @[GameLogic.scala 155:39]
  wire  _GEN_730 = kill_5_0 ? _GEN_726 : _GEN_680; // @[GameLogic.scala 155:39]
  wire  _GEN_732 = kill_5_3 & _GEN_686; // @[GameLogic.scala 157:41]
  wire  _GEN_733 = kill_5_3 ? _GEN_687 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_734 = kill_5_3 & _GEN_688; // @[GameLogic.scala 157:41]
  wire  _GEN_736 = kill_5_1 ? _GEN_732 : _GEN_686; // @[GameLogic.scala 155:39]
  wire  _GEN_737 = kill_5_1 ? _GEN_733 : _GEN_687; // @[GameLogic.scala 155:39]
  wire  _GEN_738 = kill_5_1 ? _GEN_734 : _GEN_688; // @[GameLogic.scala 155:39]
  wire  _GEN_740 = kill_5_3 & _GEN_694; // @[GameLogic.scala 157:41]
  wire  _GEN_741 = kill_5_3 ? _GEN_695 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_742 = kill_5_3 & _GEN_696; // @[GameLogic.scala 157:41]
  wire  _GEN_744 = kill_5_2 ? _GEN_740 : _GEN_694; // @[GameLogic.scala 155:39]
  wire  _GEN_745 = kill_5_2 ? _GEN_741 : _GEN_695; // @[GameLogic.scala 155:39]
  wire  _GEN_746 = kill_5_2 ? _GEN_742 : _GEN_696; // @[GameLogic.scala 155:39]
  wire  _GEN_748 = kill_5_3 & _GEN_702; // @[GameLogic.scala 157:41]
  wire  _GEN_749 = kill_5_3 ? _GEN_703 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_750 = kill_5_3 & _GEN_704; // @[GameLogic.scala 157:41]
  wire  _GEN_752 = kill_5_3 ? _GEN_748 : _GEN_702; // @[GameLogic.scala 155:39]
  wire  _GEN_753 = kill_5_3 ? _GEN_749 : _GEN_703; // @[GameLogic.scala 155:39]
  wire  _GEN_754 = kill_5_3 ? _GEN_750 : _GEN_704; // @[GameLogic.scala 155:39]
  wire  _GEN_756 = kill_5_3 & _GEN_710; // @[GameLogic.scala 157:41]
  wire  _GEN_757 = kill_5_3 ? _GEN_711 : 1'h1; // @[GameLogic.scala 157:41]
  wire  _GEN_758 = kill_5_3 & _GEN_712; // @[GameLogic.scala 157:41]
  wire  _GEN_760 = kill_5_4 ? _GEN_756 : _GEN_710; // @[GameLogic.scala 155:39]
  wire  _GEN_761 = kill_5_4 ? _GEN_757 : _GEN_711; // @[GameLogic.scala 155:39]
  wire  _GEN_762 = kill_5_4 ? _GEN_758 : _GEN_712; // @[GameLogic.scala 155:39]
  wire [10:0] _GEN_4457 = {{4{Randomizer_31_io_out[6]}},Randomizer_31_io_out}; // @[GameLogic.scala 196:51]
  wire [10:0] _T_810 = $signed(_GEN_4457) + $signed(Ystart_17); // @[GameLogic.scala 196:51]
  wire  _GEN_774 = kill_9_0 ? 1'h0 : _GEN_728; // @[GameLogic.scala 174:39]
  wire  _GEN_775 = kill_9_0 | _GEN_729; // @[GameLogic.scala 174:39]
  wire  _GEN_776 = kill_9_0 ? 1'h0 : _GEN_730; // @[GameLogic.scala 174:39]
  wire  _GEN_777 = kill_9_1 ? 1'h0 : _GEN_736; // @[GameLogic.scala 174:39]
  wire  _GEN_778 = kill_9_1 | _GEN_737; // @[GameLogic.scala 174:39]
  wire  _GEN_779 = kill_9_1 ? 1'h0 : _GEN_738; // @[GameLogic.scala 174:39]
  wire  _GEN_780 = kill_9_2 ? 1'h0 : _GEN_744; // @[GameLogic.scala 174:39]
  wire  _GEN_781 = kill_9_2 | _GEN_745; // @[GameLogic.scala 174:39]
  wire  _GEN_782 = kill_9_2 ? 1'h0 : _GEN_746; // @[GameLogic.scala 174:39]
  wire  _GEN_789 = _T_706 ? _GEN_774 : shotInteract_0; // @[GameLogic.scala 881:27]
  wire  _GEN_790 = _T_706 ? _GEN_775 : shotPop_0; // @[GameLogic.scala 881:27]
  wire  _GEN_791 = _T_706 ? _GEN_776 : spriteVisibleReg_2; // @[GameLogic.scala 881:27]
  wire  _GEN_792 = _T_706 ? _GEN_777 : shotInteract_1; // @[GameLogic.scala 881:27]
  wire  _GEN_793 = _T_706 ? _GEN_778 : shotPop_1; // @[GameLogic.scala 881:27]
  wire  _GEN_794 = _T_706 ? _GEN_779 : spriteVisibleReg_3; // @[GameLogic.scala 881:27]
  wire  _GEN_795 = _T_706 ? _GEN_780 : shotInteract_2; // @[GameLogic.scala 881:27]
  wire  _GEN_796 = _T_706 ? _GEN_781 : shotPop_2; // @[GameLogic.scala 881:27]
  wire  _GEN_797 = _T_706 ? _GEN_782 : spriteVisibleReg_4; // @[GameLogic.scala 881:27]
  wire  _GEN_798 = _T_706 ? _GEN_752 : shotInteract_3; // @[GameLogic.scala 881:27]
  wire  _GEN_799 = _T_706 ? _GEN_753 : shotPop_3; // @[GameLogic.scala 881:27]
  wire  _GEN_800 = _T_706 ? _GEN_754 : spriteVisibleReg_5; // @[GameLogic.scala 881:27]
  wire  _GEN_801 = _T_706 ? _GEN_760 : shotInteract_4; // @[GameLogic.scala 881:27]
  wire  _GEN_802 = _T_706 ? _GEN_761 : shotPop_4; // @[GameLogic.scala 881:27]
  wire  _GEN_803 = _T_706 ? _GEN_762 : spriteVisibleReg_6; // @[GameLogic.scala 881:27]
  wire  _T_815 = $signed(Ystart_17) <= 11'sh60; // @[GameLogic.scala 350:25]
  wire  _T_816 = $signed(Ystart_17) >= 11'sh120; // @[GameLogic.scala 352:31]
  wire  _GEN_824 = _T_816 | planetUp; // @[GameLogic.scala 352:43]
  wire  _GEN_825 = _T_815 ? 1'h0 : _GEN_824; // @[GameLogic.scala 350:37]
  wire  _T_817 = ~planetUp; // @[GameLogic.scala 355:44]
  wire [4:0] _T_820 = 5'sh0 - 5'sh1; // @[GameLogic.scala 355:69]
  wire [4:0] _T_821 = _T_817 ? $signed(5'sh1) : $signed(_T_820); // @[GameLogic.scala 355:43]
  wire [10:0] _GEN_4459 = {{6{_T_821[4]}},_T_821}; // @[GameLogic.scala 355:38]
  wire [10:0] _T_824 = $signed(Ystart_17) + $signed(_GEN_4459); // @[GameLogic.scala 355:38]
  wire  _T_825 = $signed(Xstart_17) > 11'sh1e0; // @[GameLogic.scala 356:42]
  wire [10:0] _T_828 = $signed(Xstart_17) - 11'sh1; // @[GameLogic.scala 356:69]
  wire  _T_830 = ~astInteract_10; // @[GameLogic.scala 363:10]
  wire  _T_833 = _T_513 & _T_688; // @[GameLogic.scala 364:26]
  wire [9:0] _T_840 = 10'sh160 - 10'sh40; // @[GameLogic.scala 368:54]
  wire  _T_841 = $signed(Randomizer_32_io_out) >= $signed(_T_840); // @[GameLogic.scala 368:45]
  wire [9:0] _T_845 = _T_841 ? $signed(_T_840) : $signed(Randomizer_32_io_out); // @[GameLogic.scala 368:30]
  wire  _GEN_826 = _T_833 | _GEN_28; // @[GameLogic.scala 364:45]
  wire  _GEN_827 = _T_833 | _GEN_29; // @[GameLogic.scala 364:45]
  wire [4:0] _T_848 = planetHp - 5'h1; // @[GameLogic.scala 378:32]
  wire [4:0] _GEN_834 = _T_688 ? _T_848 : planetHp; // @[GameLogic.scala 377:30]
  wire [4:0] _GEN_835 = kill_10_0 ? _GEN_834 : planetHp; // @[GameLogic.scala 375:36]
  wire  _GEN_836 = kill_10_0 ? 1'h0 : _GEN_789; // @[GameLogic.scala 375:36]
  wire  _GEN_837 = kill_10_0 | _GEN_790; // @[GameLogic.scala 375:36]
  wire  _GEN_838 = kill_10_0 ? 1'h0 : _GEN_791; // @[GameLogic.scala 375:36]
  wire [4:0] _GEN_839 = _T_688 ? _T_848 : _GEN_835; // @[GameLogic.scala 377:30]
  wire [4:0] _GEN_840 = kill_10_1 ? _GEN_839 : _GEN_835; // @[GameLogic.scala 375:36]
  wire  _GEN_841 = kill_10_1 ? 1'h0 : _GEN_792; // @[GameLogic.scala 375:36]
  wire  _GEN_842 = kill_10_1 | _GEN_793; // @[GameLogic.scala 375:36]
  wire  _GEN_843 = kill_10_1 ? 1'h0 : _GEN_794; // @[GameLogic.scala 375:36]
  wire  _GEN_846 = kill_10_2 ? 1'h0 : _GEN_795; // @[GameLogic.scala 375:36]
  wire  _GEN_847 = kill_10_2 | _GEN_796; // @[GameLogic.scala 375:36]
  wire  _GEN_848 = kill_10_2 ? 1'h0 : _GEN_797; // @[GameLogic.scala 375:36]
  wire  _GEN_851 = kill_10_3 ? 1'h0 : _GEN_798; // @[GameLogic.scala 375:36]
  wire  _GEN_852 = kill_10_3 | _GEN_799; // @[GameLogic.scala 375:36]
  wire  _GEN_853 = kill_10_3 ? 1'h0 : _GEN_800; // @[GameLogic.scala 375:36]
  wire  _GEN_856 = kill_10_4 ? 1'h0 : _GEN_801; // @[GameLogic.scala 375:36]
  wire  _GEN_857 = kill_10_4 | _GEN_802; // @[GameLogic.scala 375:36]
  wire  _GEN_858 = kill_10_4 ? 1'h0 : _GEN_803; // @[GameLogic.scala 375:36]
  wire  _T_862 = 4'ha == stateReg; // @[Conditional.scala 37:30]
  wire  _T_863 = hp > 4'h0; // @[GameLogic.scala 899:15]
  wire  _T_864 = $signed(Ystart_0) < 11'sh160; // @[GameLogic.scala 902:30]
  wire [10:0] _T_867 = $signed(Ystart_0) + 11'sh3; // @[GameLogic.scala 903:44]
  wire  _T_868 = $signed(Ystart_0) > 11'sh60; // @[GameLogic.scala 907:32]
  wire [10:0] _T_871 = $signed(Ystart_0) - 11'sh3; // @[GameLogic.scala 908:46]
  wire [9:0] _T_874 = 10'sh1c0 - 10'sh10; // @[GameLogic.scala 912:42]
  wire [10:0] _GEN_4461 = {{1{_T_874[9]}},_T_874}; // @[GameLogic.scala 912:30]
  wire  _T_875 = $signed(Xstart_0) < $signed(_GEN_4461); // @[GameLogic.scala 912:30]
  wire [10:0] _T_878 = $signed(Xstart_0) + 11'sh3; // @[GameLogic.scala 913:44]
  wire  _T_882 = $signed(Xstart_0) > 11'sh21; // @[GameLogic.scala 918:32]
  wire [10:0] _T_885 = $signed(Xstart_0) - 11'sh3; // @[GameLogic.scala 919:46]
  wire  _T_886 = 4'hb == stateReg; // @[Conditional.scala 37:30]
  wire [10:0] _T_889 = $signed(Xstart_2) + 11'sha; // @[GameLogic.scala 930:64]
  wire  _T_890 = $signed(Xstart_2) >= 11'sh280; // @[GameLogic.scala 266:36]
  wire  _GEN_872 = _T_890 ? 1'h0 : spriteVisibleReg_2; // @[GameLogic.scala 266:49]
  wire  _GEN_873 = _T_890 ? 1'h0 : shotInteract_0; // @[GameLogic.scala 266:49]
  wire  _GEN_874 = _T_890 | shotPop_0; // @[GameLogic.scala 266:49]
  wire [10:0] _T_893 = $signed(Xstart_3) + 11'sha; // @[GameLogic.scala 930:64]
  wire  _T_894 = $signed(Xstart_3) >= 11'sh280; // @[GameLogic.scala 266:36]
  wire  _GEN_875 = _T_894 ? 1'h0 : spriteVisibleReg_3; // @[GameLogic.scala 266:49]
  wire  _GEN_876 = _T_894 ? 1'h0 : shotInteract_1; // @[GameLogic.scala 266:49]
  wire  _GEN_877 = _T_894 | shotPop_1; // @[GameLogic.scala 266:49]
  wire [10:0] _T_897 = $signed(Xstart_4) + 11'sha; // @[GameLogic.scala 930:64]
  wire  _T_898 = $signed(Xstart_4) >= 11'sh280; // @[GameLogic.scala 266:36]
  wire  _GEN_878 = _T_898 ? 1'h0 : spriteVisibleReg_4; // @[GameLogic.scala 266:49]
  wire  _GEN_879 = _T_898 ? 1'h0 : shotInteract_2; // @[GameLogic.scala 266:49]
  wire  _GEN_880 = _T_898 | shotPop_2; // @[GameLogic.scala 266:49]
  wire [10:0] _T_901 = $signed(Xstart_5) + 11'sha; // @[GameLogic.scala 930:64]
  wire  _T_902 = $signed(Xstart_5) >= 11'sh280; // @[GameLogic.scala 266:36]
  wire  _GEN_881 = _T_902 ? 1'h0 : spriteVisibleReg_5; // @[GameLogic.scala 266:49]
  wire  _GEN_882 = _T_902 ? 1'h0 : shotInteract_3; // @[GameLogic.scala 266:49]
  wire  _GEN_883 = _T_902 | shotPop_3; // @[GameLogic.scala 266:49]
  wire [10:0] _T_905 = $signed(Xstart_6) + 11'sh1e; // @[GameLogic.scala 930:64]
  wire  _T_906 = $signed(Xstart_6) >= 11'sh280; // @[GameLogic.scala 266:36]
  wire  _GEN_884 = _T_906 ? 1'h0 : spriteVisibleReg_6; // @[GameLogic.scala 266:49]
  wire  _GEN_885 = _T_906 ? 1'h0 : shotInteract_4; // @[GameLogic.scala 266:49]
  wire  _GEN_886 = _T_906 | shotPop_4; // @[GameLogic.scala 266:49]
  wire  _T_908 = $signed(shotCntBig) > 3'sh0; // @[GameLogic.scala 934:37]
  wire  _T_909 = io_sw_1 & _T_908; // @[GameLogic.scala 934:23]
  wire  _T_911 = btnCReg & _T_908; // @[GameLogic.scala 246:18]
  wire  _GEN_887 = _T_911 | shotLoad; // @[GameLogic.scala 246:39]
  reg [10:0] _T_912; // @[GameLogic.scala 251:43]
  wire [10:0] _T_916 = $signed(_T_912) + 11'sh10; // @[GameLogic.scala 251:59]
  reg [10:0] _T_917; // @[GameLogic.scala 252:43]
  wire  _T_918 = ~btnCReg; // @[GameLogic.scala 255:22]
  wire  _T_919 = shotLoad & _T_918; // @[GameLogic.scala 255:19]
  wire [2:0] _T_922 = $signed(shotCntBig) - 3'sh1; // @[GameLogic.scala 258:32]
  wire  _GEN_890 = _T_919 | _GEN_881; // @[GameLogic.scala 255:32]
  wire  _GEN_893 = _T_919 ? 1'h0 : _GEN_883; // @[GameLogic.scala 255:32]
  wire  _GEN_894 = _T_919 | _GEN_882; // @[GameLogic.scala 255:32]
  wire  _GEN_898 = shotPop_3 ? _GEN_890 : _GEN_881; // @[GameLogic.scala 936:28]
  wire  _GEN_900 = shotPop_3 ? _GEN_893 : _GEN_883; // @[GameLogic.scala 936:28]
  wire  _GEN_901 = shotPop_3 ? _GEN_894 : _GEN_882; // @[GameLogic.scala 936:28]
  wire  _T_923 = $signed(shotCntFast) > 3'sh0; // @[GameLogic.scala 939:44]
  wire  _T_924 = io_sw_2 & _T_923; // @[GameLogic.scala 939:29]
  wire  _T_926 = btnCReg & _T_923; // @[GameLogic.scala 227:18]
  wire  _GEN_902 = _T_926 | shotLoad; // @[GameLogic.scala 227:40]
  reg [10:0] _T_927; // @[GameLogic.scala 232:43]
  wire [10:0] _T_931 = $signed(_T_927) + 11'sh10; // @[GameLogic.scala 232:59]
  reg [10:0] _T_932; // @[GameLogic.scala 233:43]
  wire [2:0] _T_937 = $signed(shotCntFast) - 3'sh1; // @[GameLogic.scala 239:34]
  wire  _GEN_905 = _T_919 | _GEN_884; // @[GameLogic.scala 236:32]
  wire  _GEN_908 = _T_919 ? 1'h0 : _GEN_886; // @[GameLogic.scala 236:32]
  wire  _GEN_909 = _T_919 | _GEN_885; // @[GameLogic.scala 236:32]
  wire  _GEN_913 = shotPop_4 ? _GEN_905 : _GEN_884; // @[GameLogic.scala 941:28]
  wire  _GEN_915 = shotPop_4 ? _GEN_908 : _GEN_886; // @[GameLogic.scala 941:28]
  wire  _GEN_916 = shotPop_4 ? _GEN_909 : _GEN_885; // @[GameLogic.scala 941:28]
  wire  _T_938 = $signed(shotCnt) > 10'sh0; // @[GameLogic.scala 206:29]
  wire  _T_939 = btnCReg & _T_938; // @[GameLogic.scala 206:18]
  wire  _GEN_917 = _T_939 | shotLoad; // @[GameLogic.scala 206:36]
  reg [10:0] _T_940; // @[GameLogic.scala 211:43]
  wire [10:0] _T_944 = $signed(_T_940) + 11'sh10; // @[GameLogic.scala 211:59]
  reg [10:0] _T_945; // @[GameLogic.scala 212:43]
  wire [9:0] _T_950 = $signed(shotCnt) - 10'sh1; // @[GameLogic.scala 218:26]
  wire  _GEN_920 = _T_919 | _GEN_872; // @[GameLogic.scala 215:32]
  wire  _GEN_923 = _T_919 ? 1'h0 : _GEN_874; // @[GameLogic.scala 215:32]
  wire  _GEN_924 = _T_919 | _GEN_873; // @[GameLogic.scala 215:32]
  wire [1:0] _GEN_925 = _T_919 ? 2'h1 : 2'h2; // @[GameLogic.scala 215:32]
  reg [10:0] _T_953; // @[GameLogic.scala 211:43]
  wire [10:0] _T_957 = $signed(_T_953) + 11'sh10; // @[GameLogic.scala 211:59]
  reg [10:0] _T_958; // @[GameLogic.scala 212:43]
  wire  _GEN_929 = _T_919 | _GEN_875; // @[GameLogic.scala 215:32]
  wire  _GEN_932 = _T_919 ? 1'h0 : _GEN_877; // @[GameLogic.scala 215:32]
  wire  _GEN_933 = _T_919 | _GEN_876; // @[GameLogic.scala 215:32]
  reg [10:0] _T_966; // @[GameLogic.scala 211:43]
  wire [10:0] _T_970 = $signed(_T_966) + 11'sh10; // @[GameLogic.scala 211:59]
  reg [10:0] _T_971; // @[GameLogic.scala 212:43]
  wire  _GEN_938 = _T_919 | _GEN_878; // @[GameLogic.scala 215:32]
  wire  _GEN_941 = _T_919 ? 1'h0 : _GEN_880; // @[GameLogic.scala 215:32]
  wire  _GEN_942 = _T_919 | _GEN_879; // @[GameLogic.scala 215:32]
  wire  _GEN_947 = shotPop_2 ? _GEN_938 : _GEN_878; // @[GameLogic.scala 950:34]
  wire  _GEN_949 = shotPop_2 ? _GEN_941 : _GEN_880; // @[GameLogic.scala 950:34]
  wire  _GEN_950 = shotPop_2 ? _GEN_942 : _GEN_879; // @[GameLogic.scala 950:34]
  wire [1:0] _GEN_951 = shotPop_2 ? _GEN_925 : 2'h2; // @[GameLogic.scala 950:34]
  wire  _GEN_955 = shotPop_1 ? _GEN_929 : _GEN_875; // @[GameLogic.scala 948:34]
  wire  _GEN_957 = shotPop_1 ? _GEN_932 : _GEN_877; // @[GameLogic.scala 948:34]
  wire  _GEN_958 = shotPop_1 ? _GEN_933 : _GEN_876; // @[GameLogic.scala 948:34]
  wire [1:0] _GEN_959 = shotPop_1 ? _GEN_925 : _GEN_951; // @[GameLogic.scala 948:34]
  wire  _GEN_962 = shotPop_1 ? _GEN_878 : _GEN_947; // @[GameLogic.scala 948:34]
  wire  _GEN_963 = shotPop_1 ? _GEN_880 : _GEN_949; // @[GameLogic.scala 948:34]
  wire  _GEN_964 = shotPop_1 ? _GEN_879 : _GEN_950; // @[GameLogic.scala 948:34]
  wire  _GEN_968 = shotPop_0 ? _GEN_920 : _GEN_872; // @[GameLogic.scala 946:28]
  wire  _GEN_970 = shotPop_0 ? _GEN_923 : _GEN_874; // @[GameLogic.scala 946:28]
  wire  _GEN_971 = shotPop_0 ? _GEN_924 : _GEN_873; // @[GameLogic.scala 946:28]
  wire [1:0] _GEN_972 = shotPop_0 ? _GEN_925 : _GEN_959; // @[GameLogic.scala 946:28]
  wire  _GEN_975 = shotPop_0 ? _GEN_875 : _GEN_955; // @[GameLogic.scala 946:28]
  wire  _GEN_976 = shotPop_0 ? _GEN_877 : _GEN_957; // @[GameLogic.scala 946:28]
  wire  _GEN_977 = shotPop_0 ? _GEN_876 : _GEN_958; // @[GameLogic.scala 946:28]
  wire  _GEN_980 = shotPop_0 ? _GEN_878 : _GEN_962; // @[GameLogic.scala 946:28]
  wire  _GEN_981 = shotPop_0 ? _GEN_880 : _GEN_963; // @[GameLogic.scala 946:28]
  wire  _GEN_982 = shotPop_0 ? _GEN_879 : _GEN_964; // @[GameLogic.scala 946:28]
  wire  _GEN_987 = _T_924 ? _GEN_913 : _GEN_884; // @[GameLogic.scala 939:51]
  wire  _GEN_989 = _T_924 ? _GEN_915 : _GEN_886; // @[GameLogic.scala 939:51]
  wire  _GEN_990 = _T_924 ? _GEN_916 : _GEN_885; // @[GameLogic.scala 939:51]
  wire  _GEN_993 = _T_924 ? _GEN_872 : _GEN_968; // @[GameLogic.scala 939:51]
  wire  _GEN_995 = _T_924 ? _GEN_874 : _GEN_970; // @[GameLogic.scala 939:51]
  wire  _GEN_996 = _T_924 ? _GEN_873 : _GEN_971; // @[GameLogic.scala 939:51]
  wire [1:0] _GEN_997 = _T_924 ? 2'h2 : _GEN_972; // @[GameLogic.scala 939:51]
  wire  _GEN_1000 = _T_924 ? _GEN_875 : _GEN_975; // @[GameLogic.scala 939:51]
  wire  _GEN_1001 = _T_924 ? _GEN_877 : _GEN_976; // @[GameLogic.scala 939:51]
  wire  _GEN_1002 = _T_924 ? _GEN_876 : _GEN_977; // @[GameLogic.scala 939:51]
  wire  _GEN_1005 = _T_924 ? _GEN_878 : _GEN_980; // @[GameLogic.scala 939:51]
  wire  _GEN_1006 = _T_924 ? _GEN_880 : _GEN_981; // @[GameLogic.scala 939:51]
  wire  _GEN_1007 = _T_924 ? _GEN_879 : _GEN_982; // @[GameLogic.scala 939:51]
  wire  _GEN_1012 = _T_909 ? _GEN_898 : _GEN_881; // @[GameLogic.scala 934:44]
  wire  _GEN_1014 = _T_909 ? _GEN_900 : _GEN_883; // @[GameLogic.scala 934:44]
  wire  _GEN_1015 = _T_909 ? _GEN_901 : _GEN_882; // @[GameLogic.scala 934:44]
  wire  _GEN_1018 = _T_909 ? _GEN_884 : _GEN_987; // @[GameLogic.scala 934:44]
  wire  _GEN_1020 = _T_909 ? _GEN_886 : _GEN_989; // @[GameLogic.scala 934:44]
  wire  _GEN_1021 = _T_909 ? _GEN_885 : _GEN_990; // @[GameLogic.scala 934:44]
  wire  _GEN_1024 = _T_909 ? _GEN_872 : _GEN_993; // @[GameLogic.scala 934:44]
  wire  _GEN_1026 = _T_909 ? _GEN_874 : _GEN_995; // @[GameLogic.scala 934:44]
  wire  _GEN_1027 = _T_909 ? _GEN_873 : _GEN_996; // @[GameLogic.scala 934:44]
  wire [1:0] _GEN_1028 = _T_909 ? 2'h2 : _GEN_997; // @[GameLogic.scala 934:44]
  wire  _GEN_1031 = _T_909 ? _GEN_875 : _GEN_1000; // @[GameLogic.scala 934:44]
  wire  _GEN_1032 = _T_909 ? _GEN_877 : _GEN_1001; // @[GameLogic.scala 934:44]
  wire  _GEN_1033 = _T_909 ? _GEN_876 : _GEN_1002; // @[GameLogic.scala 934:44]
  wire  _GEN_1036 = _T_909 ? _GEN_878 : _GEN_1005; // @[GameLogic.scala 934:44]
  wire  _GEN_1037 = _T_909 ? _GEN_880 : _GEN_1006; // @[GameLogic.scala 934:44]
  wire  _GEN_1038 = _T_909 ? _GEN_879 : _GEN_1007; // @[GameLogic.scala 934:44]
  wire  _GEN_1043 = _T_863 ? _GEN_1012 : _GEN_881; // @[GameLogic.scala 933:22]
  wire  _GEN_1045 = _T_863 ? _GEN_1014 : _GEN_883; // @[GameLogic.scala 933:22]
  wire  _GEN_1046 = _T_863 ? _GEN_1015 : _GEN_882; // @[GameLogic.scala 933:22]
  wire  _GEN_1049 = _T_863 ? _GEN_1018 : _GEN_884; // @[GameLogic.scala 933:22]
  wire  _GEN_1051 = _T_863 ? _GEN_1020 : _GEN_886; // @[GameLogic.scala 933:22]
  wire  _GEN_1052 = _T_863 ? _GEN_1021 : _GEN_885; // @[GameLogic.scala 933:22]
  wire  _GEN_1055 = _T_863 ? _GEN_1024 : _GEN_872; // @[GameLogic.scala 933:22]
  wire  _GEN_1057 = _T_863 ? _GEN_1026 : _GEN_874; // @[GameLogic.scala 933:22]
  wire  _GEN_1058 = _T_863 ? _GEN_1027 : _GEN_873; // @[GameLogic.scala 933:22]
  wire [1:0] _GEN_1059 = _T_863 ? _GEN_1028 : 2'h2; // @[GameLogic.scala 933:22]
  wire  _GEN_1062 = _T_863 ? _GEN_1031 : _GEN_875; // @[GameLogic.scala 933:22]
  wire  _GEN_1063 = _T_863 ? _GEN_1032 : _GEN_877; // @[GameLogic.scala 933:22]
  wire  _GEN_1064 = _T_863 ? _GEN_1033 : _GEN_876; // @[GameLogic.scala 933:22]
  wire  _GEN_1067 = _T_863 ? _GEN_1036 : _GEN_878; // @[GameLogic.scala 933:22]
  wire  _GEN_1068 = _T_863 ? _GEN_1037 : _GEN_880; // @[GameLogic.scala 933:22]
  wire  _GEN_1069 = _T_863 ? _GEN_1038 : _GEN_879; // @[GameLogic.scala 933:22]
  wire  _T_977 = 4'hc == stateReg; // @[Conditional.scala 37:30]
  reg  _T_978; // @[GameLogic.scala 116:23]
  reg  _T_979; // @[GameLogic.scala 117:23]
  reg [2:0] _T_980; // @[GameLogic.scala 119:25]
  reg [2:0] _T_981; // @[GameLogic.scala 120:25]
  reg [2:0] _T_982; // @[GameLogic.scala 121:25]
  wire  _T_983 = $signed(Xstart_125) > 11'sh2a0; // @[GameLogic.scala 123:26]
  wire  _T_984 = $signed(Xstart_126) > 11'sh2a0; // @[GameLogic.scala 126:26]
  wire  _T_985 = $signed(Xstart_127) > 11'sh2a0; // @[GameLogic.scala 129:26]
  wire [4:0] _GEN_4462 = {{2{_T_980[2]}},_T_980}; // @[GameLogic.scala 132:35]
  wire [4:0] _T_988 = 5'sha + $signed(_GEN_4462); // @[GameLogic.scala 132:35]
  wire [10:0] _GEN_4463 = {{6{_T_988[4]}},_T_988}; // @[GameLogic.scala 110:44]
  wire [10:0] _T_991 = $signed(Xstart_125) - $signed(_GEN_4463); // @[GameLogic.scala 110:44]
  wire  _T_992 = $signed(Xstart_125) <= 11'sh2; // @[GameLogic.scala 97:28]
  wire  _T_997 = $signed(Randomizer_35_io_out) <= 6'sh8; // @[GameLogic.scala 101:27]
  wire  _T_998 = $signed(Xstart_125) <= 11'sh160; // @[GameLogic.scala 134:26]
  wire  _GEN_1078 = _T_998 | _T_978; // @[GameLogic.scala 134:38]
  wire  _T_999 = $signed(Xstart_126) <= 11'sh160; // @[GameLogic.scala 137:26]
  wire  _GEN_1079 = _T_999 | _T_979; // @[GameLogic.scala 137:38]
  wire [4:0] _GEN_4465 = {{2{_T_981[2]}},_T_981}; // @[GameLogic.scala 141:36]
  wire [4:0] _T_1003 = 5'sh8 + $signed(_GEN_4465); // @[GameLogic.scala 141:36]
  wire [10:0] _GEN_4466 = {{6{_T_1003[4]}},_T_1003}; // @[GameLogic.scala 110:44]
  wire [10:0] _T_1006 = $signed(Xstart_126) - $signed(_GEN_4466); // @[GameLogic.scala 110:44]
  wire  _T_1007 = $signed(Xstart_126) <= 11'sh2; // @[GameLogic.scala 97:28]
  wire  _T_1012 = $signed(Randomizer_37_io_out) <= 6'sh8; // @[GameLogic.scala 101:27]
  wire [3:0] _GEN_4468 = {{1{_T_982[2]}},_T_982}; // @[GameLogic.scala 144:36]
  wire [3:0] _T_1016 = 4'sh6 + $signed(_GEN_4468); // @[GameLogic.scala 144:36]
  wire [10:0] _GEN_4469 = {{7{_T_1016[3]}},_T_1016}; // @[GameLogic.scala 110:44]
  wire [10:0] _T_1019 = $signed(Xstart_127) - $signed(_GEN_4469); // @[GameLogic.scala 110:44]
  wire  _T_1020 = $signed(Xstart_127) <= 11'sh2; // @[GameLogic.scala 97:28]
  wire  _T_1025 = $signed(Randomizer_39_io_out) <= 6'sh8; // @[GameLogic.scala 101:27]
  wire  _T_1026 = $signed(cnt) == 10'sh5; // @[GameLogic.scala 961:16]
  wire  _T_1027 = count5 == 8'h1; // @[GameLogic.scala 964:19]
  reg  _T_1028; // @[GameLogic.scala 116:23]
  reg  _T_1029; // @[GameLogic.scala 117:23]
  reg [2:0] _T_1030; // @[GameLogic.scala 119:25]
  reg [2:0] _T_1031; // @[GameLogic.scala 120:25]
  reg [2:0] _T_1032; // @[GameLogic.scala 121:25]
  wire  _T_1033 = $signed(Xstart_122) > 11'sh2a0; // @[GameLogic.scala 123:26]
  wire  _T_1034 = $signed(Xstart_123) > 11'sh2a0; // @[GameLogic.scala 126:26]
  wire  _T_1035 = $signed(Xstart_124) > 11'sh2a0; // @[GameLogic.scala 129:26]
  wire [4:0] _GEN_4471 = {{2{_T_1030[2]}},_T_1030}; // @[GameLogic.scala 132:35]
  wire [4:0] _T_1038 = 5'sha + $signed(_GEN_4471); // @[GameLogic.scala 132:35]
  wire [10:0] _GEN_4472 = {{6{_T_1038[4]}},_T_1038}; // @[GameLogic.scala 110:44]
  wire [10:0] _T_1041 = $signed(Xstart_122) - $signed(_GEN_4472); // @[GameLogic.scala 110:44]
  wire  _T_1042 = $signed(Xstart_122) <= 11'sh2; // @[GameLogic.scala 97:28]
  wire  _T_1047 = $signed(Randomizer_42_io_out) <= 6'sh8; // @[GameLogic.scala 101:27]
  wire  _T_1048 = $signed(Xstart_122) <= 11'sh160; // @[GameLogic.scala 134:26]
  wire  _GEN_1107 = _T_1048 | _T_1028; // @[GameLogic.scala 134:38]
  wire  _T_1049 = $signed(Xstart_123) <= 11'sh160; // @[GameLogic.scala 137:26]
  wire  _GEN_1108 = _T_1049 | _T_1029; // @[GameLogic.scala 137:38]
  wire [4:0] _GEN_4474 = {{2{_T_1031[2]}},_T_1031}; // @[GameLogic.scala 141:36]
  wire [4:0] _T_1053 = 5'sh8 + $signed(_GEN_4474); // @[GameLogic.scala 141:36]
  wire [10:0] _GEN_4475 = {{6{_T_1053[4]}},_T_1053}; // @[GameLogic.scala 110:44]
  wire [10:0] _T_1056 = $signed(Xstart_123) - $signed(_GEN_4475); // @[GameLogic.scala 110:44]
  wire  _T_1057 = $signed(Xstart_123) <= 11'sh2; // @[GameLogic.scala 97:28]
  wire  _T_1062 = $signed(Randomizer_44_io_out) <= 6'sh8; // @[GameLogic.scala 101:27]
  wire [3:0] _GEN_4477 = {{1{_T_1032[2]}},_T_1032}; // @[GameLogic.scala 144:36]
  wire [3:0] _T_1066 = 4'sh6 + $signed(_GEN_4477); // @[GameLogic.scala 144:36]
  wire [10:0] _GEN_4478 = {{7{_T_1066[3]}},_T_1066}; // @[GameLogic.scala 110:44]
  wire [10:0] _T_1069 = $signed(Xstart_124) - $signed(_GEN_4478); // @[GameLogic.scala 110:44]
  wire  _T_1070 = $signed(Xstart_124) <= 11'sh2; // @[GameLogic.scala 97:28]
  wire  _T_1075 = $signed(Randomizer_46_io_out) <= 6'sh8; // @[GameLogic.scala 101:27]
  wire  _T_1076 = io_btnC | io_btnL; // @[GameLogic.scala 968:28]
  wire  _T_1077 = _T_1076 | io_btnD; // @[GameLogic.scala 968:39]
  wire  _T_1078 = _T_1077 | io_btnU; // @[GameLogic.scala 968:50]
  wire  _T_1079 = _T_1078 | io_btnR; // @[GameLogic.scala 968:61]
  wire  _T_1080 = _T_1079 | start; // @[GameLogic.scala 968:19]
  wire  _T_1082 = $signed(secCnt) <= 8'sh9; // @[GameLogic.scala 969:36]
  wire  _T_1083 = _T_513 & _T_1082; // @[GameLogic.scala 969:26]
  wire  _T_1084 = level == 3'h4; // @[GameLogic.scala 969:52]
  wire  _T_1085 = _T_1083 & _T_1084; // @[GameLogic.scala 969:43]
  wire  _T_1087 = $signed(cnt) == 10'sh3c; // @[GameLogic.scala 980:16]
  wire  _T_1088 = _T_1087 & start; // @[GameLogic.scala 980:25]
  wire [7:0] _T_1091 = $signed(secCnt) + 8'sh1; // @[GameLogic.scala 981:26]
  wire  _T_1092 = $signed(secCnt) == 8'shf; // @[GameLogic.scala 982:35]
  wire  _T_1093 = io_sw_7 & _T_1092; // @[GameLogic.scala 982:25]
  wire  _T_1094 = $signed(secCnt) == 8'sh3c; // @[GameLogic.scala 982:55]
  wire  _T_1095 = _T_1093 | _T_1094; // @[GameLogic.scala 982:45]
  wire  _T_1097 = _T_1095 & _T_863; // @[GameLogic.scala 982:65]
  wire  _T_1099 = _T_1097 & _T_506; // @[GameLogic.scala 982:77]
  wire [2:0] _T_1101 = level + 3'h1; // @[GameLogic.scala 984:26]
  wire  _T_1104 = _T_1094 & _T_1084; // @[GameLogic.scala 987:36]
  wire [3:0] _GEN_1161 = _T_1099 ? 4'h3 : hp; // @[GameLogic.scala 982:93]
  wire  _GEN_1167 = _T_1099 | levelCng; // @[GameLogic.scala 982:93]
  wire [3:0] _GEN_1169 = _T_1088 ? _GEN_1161 : hp; // @[GameLogic.scala 980:35]
  wire [9:0] _T_1108 = $signed(cnt) + 10'sh1; // @[GameLogic.scala 992:41]
  wire  _T_1111 = cng ? _T_26 : show; // @[GameLogic.scala 993:18]
  wire  _T_1112 = $signed(cnt) < 10'sh7; // @[GameLogic.scala 994:21]
  wire  _T_1113 = $signed(cnt) > 10'sh1e; // @[GameLogic.scala 994:35]
  wire  _T_1114 = $signed(cnt) < 10'sh25; // @[GameLogic.scala 994:49]
  wire  _T_1115 = _T_1113 & _T_1114; // @[GameLogic.scala 994:42]
  wire  _T_1116 = _T_1112 | _T_1115; // @[GameLogic.scala 994:27]
  wire  _T_1118 = cng & _T_281; // @[GameLogic.scala 995:16]
  wire [3:0] _T_1120 = cngCnt + 4'h1; // @[GameLogic.scala 996:26]
  wire  _T_1121 = cngCnt >= 4'h5; // @[GameLogic.scala 997:21]
  wire  _T_1122 = astInteract_0 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1123 = _T_1122 & boxDetection_io_overlap_0_7; // @[GameLogic.scala 1003:50]
  wire  _T_1124 = astInteract_0 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1125 = _T_1124 & boxDetection_io_overlap_2_7; // @[GameLogic.scala 1005:59]
  wire  _T_1126 = astInteract_0 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1127 = _T_1126 & boxDetection_io_overlap_3_7; // @[GameLogic.scala 1005:59]
  wire  _T_1128 = astInteract_0 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1129 = _T_1128 & boxDetection_io_overlap_4_7; // @[GameLogic.scala 1005:59]
  wire  _T_1130 = astInteract_0 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1131 = _T_1130 & boxDetection_io_overlap_5_7; // @[GameLogic.scala 1005:59]
  wire  _T_1132 = astInteract_0 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1133 = _T_1132 & boxDetection_io_overlap_6_7; // @[GameLogic.scala 1005:59]
  wire  _T_1134 = hp > 4'h1; // @[GameLogic.scala 280:15]
  wire [10:0] _GEN_1177 = _T_1134 ? $signed(11'sh40) : $signed(Xstart_0); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1178 = _T_1134 ? $signed(11'she0) : $signed(Ystart_0); // @[GameLogic.scala 280:22]
  wire  _T_1136 = shipInteract & _T_863; // @[GameLogic.scala 285:25]
  wire [3:0] _T_1138 = hp - 4'h1; // @[GameLogic.scala 286:18]
  wire [3:0] _GEN_1179 = _T_1136 ? _T_1138 : _GEN_1169; // @[GameLogic.scala 285:38]
  wire  _GEN_1181 = _T_1136 ? 1'h0 : shipInteract; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1182 = die_0 ? $signed(_GEN_1177) : $signed(Xstart_0); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1183 = die_0 ? $signed(_GEN_1178) : $signed(Ystart_0); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1184 = die_0 ? _GEN_1179 : _GEN_1169; // @[GameLogic.scala 274:18]
  wire  _GEN_1186 = die_0 ? _GEN_1181 : shipInteract; // @[GameLogic.scala 274:18]
  wire  _T_1139 = astInteract_1 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1140 = _T_1139 & boxDetection_io_overlap_0_8; // @[GameLogic.scala 1003:50]
  wire  _T_1141 = astInteract_1 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1142 = _T_1141 & boxDetection_io_overlap_2_8; // @[GameLogic.scala 1005:59]
  wire  _T_1143 = astInteract_1 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1144 = _T_1143 & boxDetection_io_overlap_3_8; // @[GameLogic.scala 1005:59]
  wire  _T_1145 = astInteract_1 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1146 = _T_1145 & boxDetection_io_overlap_4_8; // @[GameLogic.scala 1005:59]
  wire  _T_1147 = astInteract_1 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1148 = _T_1147 & boxDetection_io_overlap_5_8; // @[GameLogic.scala 1005:59]
  wire  _T_1149 = astInteract_1 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1150 = _T_1149 & boxDetection_io_overlap_6_8; // @[GameLogic.scala 1005:59]
  wire [10:0] _GEN_1187 = _T_1134 ? $signed(11'sh40) : $signed(_GEN_1182); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1188 = _T_1134 ? $signed(11'she0) : $signed(_GEN_1183); // @[GameLogic.scala 280:22]
  wire [3:0] _GEN_1189 = _T_1136 ? _T_1138 : _GEN_1184; // @[GameLogic.scala 285:38]
  wire  _GEN_1191 = _T_1136 ? 1'h0 : _GEN_1186; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1192 = die_1 ? $signed(_GEN_1187) : $signed(_GEN_1182); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1193 = die_1 ? $signed(_GEN_1188) : $signed(_GEN_1183); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1194 = die_1 ? _GEN_1189 : _GEN_1184; // @[GameLogic.scala 274:18]
  wire  _GEN_1196 = die_1 ? _GEN_1191 : _GEN_1186; // @[GameLogic.scala 274:18]
  wire  _T_1156 = astInteract_2 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1157 = _T_1156 & boxDetection_io_overlap_0_9; // @[GameLogic.scala 1003:50]
  wire  _T_1158 = astInteract_2 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1159 = _T_1158 & boxDetection_io_overlap_2_9; // @[GameLogic.scala 1005:59]
  wire  _T_1160 = astInteract_2 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1161 = _T_1160 & boxDetection_io_overlap_3_9; // @[GameLogic.scala 1005:59]
  wire  _T_1162 = astInteract_2 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1163 = _T_1162 & boxDetection_io_overlap_4_9; // @[GameLogic.scala 1005:59]
  wire  _T_1164 = astInteract_2 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1165 = _T_1164 & boxDetection_io_overlap_5_9; // @[GameLogic.scala 1005:59]
  wire  _T_1166 = astInteract_2 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1167 = _T_1166 & boxDetection_io_overlap_6_9; // @[GameLogic.scala 1005:59]
  wire [10:0] _GEN_1197 = _T_1134 ? $signed(11'sh40) : $signed(_GEN_1192); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1198 = _T_1134 ? $signed(11'she0) : $signed(_GEN_1193); // @[GameLogic.scala 280:22]
  wire [3:0] _GEN_1199 = _T_1136 ? _T_1138 : _GEN_1194; // @[GameLogic.scala 285:38]
  wire  _GEN_1201 = _T_1136 ? 1'h0 : _GEN_1196; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1202 = die_2 ? $signed(_GEN_1197) : $signed(_GEN_1192); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1203 = die_2 ? $signed(_GEN_1198) : $signed(_GEN_1193); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1204 = die_2 ? _GEN_1199 : _GEN_1194; // @[GameLogic.scala 274:18]
  wire  _GEN_1206 = die_2 ? _GEN_1201 : _GEN_1196; // @[GameLogic.scala 274:18]
  wire  _T_1173 = astInteract_3 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1174 = _T_1173 & boxDetection_io_overlap_0_10; // @[GameLogic.scala 1003:50]
  wire  _T_1175 = astInteract_3 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1176 = _T_1175 & boxDetection_io_overlap_2_10; // @[GameLogic.scala 1005:59]
  wire  _T_1177 = astInteract_3 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1178 = _T_1177 & boxDetection_io_overlap_3_10; // @[GameLogic.scala 1005:59]
  wire  _T_1179 = astInteract_3 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1180 = _T_1179 & boxDetection_io_overlap_4_10; // @[GameLogic.scala 1005:59]
  wire  _T_1181 = astInteract_3 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1182 = _T_1181 & boxDetection_io_overlap_5_10; // @[GameLogic.scala 1005:59]
  wire  _T_1183 = astInteract_3 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1184 = _T_1183 & boxDetection_io_overlap_6_10; // @[GameLogic.scala 1005:59]
  wire [10:0] _GEN_1207 = _T_1134 ? $signed(11'sh40) : $signed(_GEN_1202); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1208 = _T_1134 ? $signed(11'she0) : $signed(_GEN_1203); // @[GameLogic.scala 280:22]
  wire [3:0] _GEN_1209 = _T_1136 ? _T_1138 : _GEN_1204; // @[GameLogic.scala 285:38]
  wire  _GEN_1211 = _T_1136 ? 1'h0 : _GEN_1206; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1212 = die_3 ? $signed(_GEN_1207) : $signed(_GEN_1202); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1213 = die_3 ? $signed(_GEN_1208) : $signed(_GEN_1203); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1214 = die_3 ? _GEN_1209 : _GEN_1204; // @[GameLogic.scala 274:18]
  wire  _GEN_1216 = die_3 ? _GEN_1211 : _GEN_1206; // @[GameLogic.scala 274:18]
  wire  _T_1190 = astInteract_4 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1191 = _T_1190 & boxDetection_io_overlap_0_11; // @[GameLogic.scala 1003:50]
  wire  _T_1192 = astInteract_4 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1193 = _T_1192 & boxDetection_io_overlap_2_11; // @[GameLogic.scala 1005:59]
  wire  _T_1194 = astInteract_4 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1195 = _T_1194 & boxDetection_io_overlap_3_11; // @[GameLogic.scala 1005:59]
  wire  _T_1196 = astInteract_4 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1197 = _T_1196 & boxDetection_io_overlap_4_11; // @[GameLogic.scala 1005:59]
  wire  _T_1198 = astInteract_4 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1199 = _T_1198 & boxDetection_io_overlap_5_11; // @[GameLogic.scala 1005:59]
  wire  _T_1200 = astInteract_4 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1201 = _T_1200 & boxDetection_io_overlap_6_11; // @[GameLogic.scala 1005:59]
  wire [10:0] _GEN_1217 = _T_1134 ? $signed(11'sh40) : $signed(_GEN_1212); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1218 = _T_1134 ? $signed(11'she0) : $signed(_GEN_1213); // @[GameLogic.scala 280:22]
  wire [3:0] _GEN_1219 = _T_1136 ? _T_1138 : _GEN_1214; // @[GameLogic.scala 285:38]
  wire  _GEN_1221 = _T_1136 ? 1'h0 : _GEN_1216; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1222 = die_4 ? $signed(_GEN_1217) : $signed(_GEN_1212); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1223 = die_4 ? $signed(_GEN_1218) : $signed(_GEN_1213); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1224 = die_4 ? _GEN_1219 : _GEN_1214; // @[GameLogic.scala 274:18]
  wire  _GEN_1226 = die_4 ? _GEN_1221 : _GEN_1216; // @[GameLogic.scala 274:18]
  wire  _T_1207 = astInteract_5 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1208 = _T_1207 & boxDetection_io_overlap_0_12; // @[GameLogic.scala 1003:50]
  wire  _T_1209 = astInteract_5 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1210 = _T_1209 & boxDetection_io_overlap_2_12; // @[GameLogic.scala 1005:59]
  wire  _T_1211 = astInteract_5 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1212 = _T_1211 & boxDetection_io_overlap_3_12; // @[GameLogic.scala 1005:59]
  wire  _T_1213 = astInteract_5 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1214 = _T_1213 & boxDetection_io_overlap_4_12; // @[GameLogic.scala 1005:59]
  wire  _T_1215 = astInteract_5 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1216 = _T_1215 & boxDetection_io_overlap_5_12; // @[GameLogic.scala 1005:59]
  wire  _T_1217 = astInteract_5 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1218 = _T_1217 & boxDetection_io_overlap_6_12; // @[GameLogic.scala 1005:59]
  wire [10:0] _GEN_1227 = _T_1134 ? $signed(11'sh40) : $signed(_GEN_1222); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1228 = _T_1134 ? $signed(11'she0) : $signed(_GEN_1223); // @[GameLogic.scala 280:22]
  wire [3:0] _GEN_1229 = _T_1136 ? _T_1138 : _GEN_1224; // @[GameLogic.scala 285:38]
  wire  _GEN_1231 = _T_1136 ? 1'h0 : _GEN_1226; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1232 = die_5 ? $signed(_GEN_1227) : $signed(_GEN_1222); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1233 = die_5 ? $signed(_GEN_1228) : $signed(_GEN_1223); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1234 = die_5 ? _GEN_1229 : _GEN_1224; // @[GameLogic.scala 274:18]
  wire  _GEN_1236 = die_5 ? _GEN_1231 : _GEN_1226; // @[GameLogic.scala 274:18]
  wire  _T_1224 = astInteract_6 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1225 = _T_1224 & boxDetection_io_overlap_0_13; // @[GameLogic.scala 1003:50]
  wire  _T_1226 = astInteract_6 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1227 = _T_1226 & boxDetection_io_overlap_2_13; // @[GameLogic.scala 1005:59]
  wire  _T_1228 = astInteract_6 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1229 = _T_1228 & boxDetection_io_overlap_3_13; // @[GameLogic.scala 1005:59]
  wire  _T_1230 = astInteract_6 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1231 = _T_1230 & boxDetection_io_overlap_4_13; // @[GameLogic.scala 1005:59]
  wire  _T_1232 = astInteract_6 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1233 = _T_1232 & boxDetection_io_overlap_5_13; // @[GameLogic.scala 1005:59]
  wire  _T_1234 = astInteract_6 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1235 = _T_1234 & boxDetection_io_overlap_6_13; // @[GameLogic.scala 1005:59]
  wire [10:0] _GEN_1237 = _T_1134 ? $signed(11'sh40) : $signed(_GEN_1232); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1238 = _T_1134 ? $signed(11'she0) : $signed(_GEN_1233); // @[GameLogic.scala 280:22]
  wire [3:0] _GEN_1239 = _T_1136 ? _T_1138 : _GEN_1234; // @[GameLogic.scala 285:38]
  wire  _GEN_1241 = _T_1136 ? 1'h0 : _GEN_1236; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1242 = die_6 ? $signed(_GEN_1237) : $signed(_GEN_1232); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1243 = die_6 ? $signed(_GEN_1238) : $signed(_GEN_1233); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1244 = die_6 ? _GEN_1239 : _GEN_1234; // @[GameLogic.scala 274:18]
  wire  _GEN_1246 = die_6 ? _GEN_1241 : _GEN_1236; // @[GameLogic.scala 274:18]
  wire  _T_1241 = astInteract_7 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1242 = _T_1241 & boxDetection_io_overlap_0_14; // @[GameLogic.scala 1003:50]
  wire  _T_1243 = astInteract_7 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1244 = _T_1243 & boxDetection_io_overlap_2_14; // @[GameLogic.scala 1005:59]
  wire  _T_1245 = astInteract_7 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1246 = _T_1245 & boxDetection_io_overlap_3_14; // @[GameLogic.scala 1005:59]
  wire  _T_1247 = astInteract_7 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1248 = _T_1247 & boxDetection_io_overlap_4_14; // @[GameLogic.scala 1005:59]
  wire  _T_1249 = astInteract_7 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1250 = _T_1249 & boxDetection_io_overlap_5_14; // @[GameLogic.scala 1005:59]
  wire  _T_1251 = astInteract_7 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1252 = _T_1251 & boxDetection_io_overlap_6_14; // @[GameLogic.scala 1005:59]
  wire [10:0] _GEN_1247 = _T_1134 ? $signed(11'sh40) : $signed(_GEN_1242); // @[GameLogic.scala 280:22]
  wire [10:0] _GEN_1248 = _T_1134 ? $signed(11'she0) : $signed(_GEN_1243); // @[GameLogic.scala 280:22]
  wire [3:0] _GEN_1249 = _T_1136 ? _T_1138 : _GEN_1244; // @[GameLogic.scala 285:38]
  wire  _GEN_1251 = _T_1136 ? 1'h0 : _GEN_1246; // @[GameLogic.scala 285:38]
  wire [10:0] _GEN_1252 = die_7 ? $signed(_GEN_1247) : $signed(_GEN_1242); // @[GameLogic.scala 274:18]
  wire [10:0] _GEN_1253 = die_7 ? $signed(_GEN_1248) : $signed(_GEN_1243); // @[GameLogic.scala 274:18]
  wire [3:0] _GEN_1254 = die_7 ? _GEN_1249 : _GEN_1244; // @[GameLogic.scala 274:18]
  wire  _GEN_1256 = die_7 ? _GEN_1251 : _GEN_1246; // @[GameLogic.scala 274:18]
  wire  _T_1258 = astInteract_8 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1259 = _T_1258 & boxDetection_io_overlap_0_15; // @[GameLogic.scala 1003:50]
  wire  _T_1260 = astInteract_8 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1261 = _T_1260 & boxDetection_io_overlap_2_15; // @[GameLogic.scala 1005:59]
  wire  _T_1262 = astInteract_8 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1263 = _T_1262 & boxDetection_io_overlap_3_15; // @[GameLogic.scala 1005:59]
  wire  _T_1264 = astInteract_8 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1265 = _T_1264 & boxDetection_io_overlap_4_15; // @[GameLogic.scala 1005:59]
  wire  _T_1266 = astInteract_8 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1267 = _T_1266 & boxDetection_io_overlap_5_15; // @[GameLogic.scala 1005:59]
  wire  _T_1268 = astInteract_8 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1269 = _T_1268 & boxDetection_io_overlap_6_15; // @[GameLogic.scala 1005:59]
  wire  _GEN_1261 = _T_1136 ? 1'h0 : _GEN_1256; // @[GameLogic.scala 285:38]
  wire  _GEN_1266 = die_8 ? _GEN_1261 : _GEN_1256; // @[GameLogic.scala 274:18]
  wire  _T_1275 = astInteract_9 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1276 = _T_1275 & boxDetection_io_overlap_0_16; // @[GameLogic.scala 1003:50]
  wire  _T_1277 = astInteract_9 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1278 = _T_1277 & boxDetection_io_overlap_2_16; // @[GameLogic.scala 1005:59]
  wire  _T_1279 = astInteract_9 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1280 = _T_1279 & boxDetection_io_overlap_3_16; // @[GameLogic.scala 1005:59]
  wire  _T_1281 = astInteract_9 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1282 = _T_1281 & boxDetection_io_overlap_4_16; // @[GameLogic.scala 1005:59]
  wire  _T_1283 = astInteract_9 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1284 = _T_1283 & boxDetection_io_overlap_5_16; // @[GameLogic.scala 1005:59]
  wire  _GEN_1271 = _T_1136 ? 1'h0 : _GEN_1266; // @[GameLogic.scala 285:38]
  wire  _GEN_1276 = die_9 ? _GEN_1271 : _GEN_1266; // @[GameLogic.scala 274:18]
  wire  _T_1292 = astInteract_10 & shipInteract; // @[GameLogic.scala 1003:34]
  wire  _T_1293 = _T_1292 & boxDetection_io_overlap_0_17; // @[GameLogic.scala 1003:50]
  wire  _T_1294 = astInteract_10 & shotInteract_0; // @[GameLogic.scala 1005:40]
  wire  _T_1295 = _T_1294 & boxDetection_io_overlap_2_17; // @[GameLogic.scala 1005:59]
  wire  _T_1296 = astInteract_10 & shotInteract_1; // @[GameLogic.scala 1005:40]
  wire  _T_1297 = _T_1296 & boxDetection_io_overlap_3_17; // @[GameLogic.scala 1005:59]
  wire  _T_1298 = astInteract_10 & shotInteract_2; // @[GameLogic.scala 1005:40]
  wire  _T_1299 = _T_1298 & boxDetection_io_overlap_4_17; // @[GameLogic.scala 1005:59]
  wire  _T_1300 = astInteract_10 & shotInteract_3; // @[GameLogic.scala 1005:40]
  wire  _T_1301 = _T_1300 & boxDetection_io_overlap_5_17; // @[GameLogic.scala 1005:59]
  wire  _T_1302 = astInteract_10 & shotInteract_4; // @[GameLogic.scala 1005:40]
  wire  _T_1303 = _T_1302 & boxDetection_io_overlap_6_17; // @[GameLogic.scala 1005:59]
  wire  _GEN_1281 = _T_1136 ? 1'h0 : _GEN_1276; // @[GameLogic.scala 285:38]
  wire  _GEN_1286 = die_10 ? _GEN_1281 : _GEN_1276; // @[GameLogic.scala 274:18]
  wire  _T_1310 = cng & _T_27; // @[GameLogic.scala 1009:16]
  wire [5:0] _T_1313 = $signed(spwnProt) + 6'sh1; // @[GameLogic.scala 1010:30]
  wire  _T_1314 = $signed(spwnProt) >= 6'sh6; // @[GameLogic.scala 1012:21]
  wire  _GEN_1288 = _T_1314 | _GEN_1286; // @[GameLogic.scala 1012:29]
  wire  _GEN_1294 = io_sw_0 | _T_1080; // @[GameLogic.scala 1016:22]
  wire  _T_1359 = $signed(shotCntFast) > 3'sh1; // @[GameLogic.scala 315:47]
  wire  _T_1360 = $signed(shotCntBig) > 3'sh1; // @[GameLogic.scala 316:46]
  wire  _T_1361 = $signed(shotCnt) > 10'sh5; // @[GameLogic.scala 317:43]
  wire  _T_1363 = $signed(shotCntFast) > 3'sh2; // @[GameLogic.scala 315:47]
  wire  _T_1364 = $signed(shotCntBig) > 3'sh2; // @[GameLogic.scala 316:46]
  wire  _T_1365 = $signed(shotCnt) > 10'sha; // @[GameLogic.scala 317:43]
  wire  _T_1366 = hp > 4'h2; // @[GameLogic.scala 318:38]
  wire [5:0] _T_1367 = 5'sh8 * 5'sh0; // @[GameLogic.scala 323:55]
  wire [6:0] _T_1368 = {{1{_T_1367[5]}},_T_1367}; // @[GameLogic.scala 323:48]
  wire [5:0] _T_1370 = _T_1368[5:0]; // @[GameLogic.scala 323:48]
  wire [7:0] _GEN_4480 = {{2{_T_1370[5]}},_T_1370}; // @[GameLogic.scala 323:42]
  wire  _T_1371 = $signed(secCnt) > $signed(_GEN_4480); // @[GameLogic.scala 323:42]
  wire [5:0] _T_1375 = 6'sh8 + $signed(_T_1367); // @[GameLogic.scala 323:79]
  wire [7:0] _GEN_4481 = {{2{_T_1375[5]}},_T_1375}; // @[GameLogic.scala 323:72]
  wire  _T_1376 = $signed(secCnt) <= $signed(_GEN_4481); // @[GameLogic.scala 323:72]
  wire  _T_1377 = _T_1371 & _T_1376; // @[GameLogic.scala 323:62]
  wire [6:0] _T_1378 = 5'sh8 * 5'sh1; // @[GameLogic.scala 323:55]
  wire [7:0] _T_1379 = {{1{_T_1378[6]}},_T_1378}; // @[GameLogic.scala 323:48]
  wire [6:0] _T_1381 = _T_1379[6:0]; // @[GameLogic.scala 323:48]
  wire [7:0] _GEN_4482 = {{1{_T_1381[6]}},_T_1381}; // @[GameLogic.scala 323:42]
  wire  _T_1382 = $signed(secCnt) > $signed(_GEN_4482); // @[GameLogic.scala 323:42]
  wire [6:0] _T_1386 = 7'sh8 + $signed(_T_1378); // @[GameLogic.scala 323:79]
  wire [7:0] _GEN_4483 = {{1{_T_1386[6]}},_T_1386}; // @[GameLogic.scala 323:72]
  wire  _T_1387 = $signed(secCnt) <= $signed(_GEN_4483); // @[GameLogic.scala 323:72]
  wire  _T_1388 = _T_1382 & _T_1387; // @[GameLogic.scala 323:62]
  wire [7:0] _T_1389 = 5'sh8 * 5'sh2; // @[GameLogic.scala 323:55]
  wire [8:0] _T_1390 = {{1{_T_1389[7]}},_T_1389}; // @[GameLogic.scala 323:48]
  wire [7:0] _T_1392 = _T_1390[7:0]; // @[GameLogic.scala 323:48]
  wire  _T_1393 = $signed(secCnt) > $signed(_T_1392); // @[GameLogic.scala 323:42]
  wire [7:0] _T_1397 = 8'sh8 + $signed(_T_1389); // @[GameLogic.scala 323:79]
  wire  _T_1398 = $signed(secCnt) <= $signed(_T_1397); // @[GameLogic.scala 323:72]
  wire  _T_1399 = _T_1393 & _T_1398; // @[GameLogic.scala 323:62]
  wire [7:0] _T_1400 = 5'sh8 * 5'sh3; // @[GameLogic.scala 323:55]
  wire [8:0] _T_1401 = {{1{_T_1400[7]}},_T_1400}; // @[GameLogic.scala 323:48]
  wire [7:0] _T_1403 = _T_1401[7:0]; // @[GameLogic.scala 323:48]
  wire  _T_1404 = $signed(secCnt) > $signed(_T_1403); // @[GameLogic.scala 323:42]
  wire [7:0] _T_1408 = 8'sh8 + $signed(_T_1400); // @[GameLogic.scala 323:79]
  wire  _T_1409 = $signed(secCnt) <= $signed(_T_1408); // @[GameLogic.scala 323:72]
  wire  _T_1410 = _T_1404 & _T_1409; // @[GameLogic.scala 323:62]
  wire [8:0] _T_1411 = 5'sh8 * 5'sh4; // @[GameLogic.scala 323:55]
  wire [9:0] _T_1412 = {{1{_T_1411[8]}},_T_1411}; // @[GameLogic.scala 323:48]
  wire [8:0] _T_1414 = _T_1412[8:0]; // @[GameLogic.scala 323:48]
  wire [8:0] _GEN_4484 = {{1{secCnt[7]}},secCnt}; // @[GameLogic.scala 323:42]
  wire  _T_1415 = $signed(_GEN_4484) > $signed(_T_1414); // @[GameLogic.scala 323:42]
  wire [8:0] _T_1419 = 9'sh8 + $signed(_T_1411); // @[GameLogic.scala 323:79]
  wire  _T_1420 = $signed(_GEN_4484) <= $signed(_T_1419); // @[GameLogic.scala 323:72]
  wire  _T_1421 = _T_1415 & _T_1420; // @[GameLogic.scala 323:62]
  wire [8:0] _T_1422 = 5'sh8 * 5'sh5; // @[GameLogic.scala 323:55]
  wire [9:0] _T_1423 = {{1{_T_1422[8]}},_T_1422}; // @[GameLogic.scala 323:48]
  wire [8:0] _T_1425 = _T_1423[8:0]; // @[GameLogic.scala 323:48]
  wire  _T_1426 = $signed(_GEN_4484) > $signed(_T_1425); // @[GameLogic.scala 323:42]
  wire [8:0] _T_1430 = 9'sh8 + $signed(_T_1422); // @[GameLogic.scala 323:79]
  wire  _T_1431 = $signed(_GEN_4484) <= $signed(_T_1430); // @[GameLogic.scala 323:72]
  wire  _T_1432 = _T_1426 & _T_1431; // @[GameLogic.scala 323:62]
  wire [8:0] _T_1433 = 5'sh8 * 5'sh6; // @[GameLogic.scala 323:55]
  wire [9:0] _T_1434 = {{1{_T_1433[8]}},_T_1433}; // @[GameLogic.scala 323:48]
  wire [8:0] _T_1436 = _T_1434[8:0]; // @[GameLogic.scala 323:48]
  wire  _T_1437 = $signed(_GEN_4484) > $signed(_T_1436); // @[GameLogic.scala 323:42]
  wire [8:0] _T_1441 = 9'sh8 + $signed(_T_1433); // @[GameLogic.scala 323:79]
  wire  _T_1442 = $signed(_GEN_4484) <= $signed(_T_1441); // @[GameLogic.scala 323:72]
  wire  _T_1443 = _T_1437 & _T_1442; // @[GameLogic.scala 323:62]
  wire [8:0] _T_1444 = 5'sh8 * 5'sh7; // @[GameLogic.scala 323:55]
  wire [9:0] _T_1445 = {{1{_T_1444[8]}},_T_1444}; // @[GameLogic.scala 323:48]
  wire [8:0] _T_1447 = _T_1445[8:0]; // @[GameLogic.scala 323:48]
  wire  _T_1448 = $signed(_GEN_4484) > $signed(_T_1447); // @[GameLogic.scala 323:42]
  wire [8:0] _T_1452 = 9'sh8 + $signed(_T_1444); // @[GameLogic.scala 323:79]
  wire  _T_1453 = $signed(_GEN_4484) <= $signed(_T_1452); // @[GameLogic.scala 323:72]
  wire  _T_1454 = _T_1448 & _T_1453; // @[GameLogic.scala 323:62]
  wire  _T_1455 = 4'hd == stateReg; // @[Conditional.scala 37:30]
  wire  _GEN_1352 = _T_977 ? _T_1111 : show; // @[Conditional.scala 39:67]
  wire  _GEN_1363 = _T_977 ? _GEN_1288 : shipInteract; // @[Conditional.scala 39:67]
  wire  _GEN_1427 = _T_977 ? _T_281 : spriteVisibleReg_26; // @[Conditional.scala 39:67]
  wire  _GEN_1430 = _T_977 ? _T_500 : spriteVisibleReg_30; // @[Conditional.scala 39:67]
  wire  _GEN_1433 = _T_977 ? _T_281 : spriteVisibleReg_27; // @[Conditional.scala 39:67]
  wire  _GEN_1436 = _T_977 ? _T_500 : spriteVisibleReg_31; // @[Conditional.scala 39:67]
  wire  _GEN_1439 = _T_977 ? _T_281 : spriteVisibleReg_28; // @[Conditional.scala 39:67]
  wire  _GEN_1442 = _T_977 ? _T_500 : spriteVisibleReg_32; // @[Conditional.scala 39:67]
  wire  _GEN_1445 = _T_977 ? _T_281 : spriteVisibleReg_29; // @[Conditional.scala 39:67]
  wire  _GEN_1448 = _T_977 ? _T_500 : spriteVisibleReg_33; // @[Conditional.scala 39:67]
  wire  _GEN_1451 = _T_977 ? _T_923 : spriteVisibleReg_72; // @[Conditional.scala 39:67]
  wire  _GEN_1452 = _T_977 ? _T_908 : spriteVisibleReg_66; // @[Conditional.scala 39:67]
  wire  _GEN_1453 = _T_977 ? _T_938 : spriteVisibleReg_57; // @[Conditional.scala 39:67]
  wire  _GEN_1454 = _T_977 ? _T_863 : spriteVisibleReg_61; // @[Conditional.scala 39:67]
  wire  _GEN_1455 = _T_977 ? _T_1359 : spriteVisibleReg_71; // @[Conditional.scala 39:67]
  wire  _GEN_1456 = _T_977 ? _T_1360 : spriteVisibleReg_65; // @[Conditional.scala 39:67]
  wire  _GEN_1457 = _T_977 ? _T_1361 : spriteVisibleReg_56; // @[Conditional.scala 39:67]
  wire  _GEN_1458 = _T_977 ? _T_1134 : spriteVisibleReg_62; // @[Conditional.scala 39:67]
  wire  _GEN_1459 = _T_977 ? _T_1363 : spriteVisibleReg_70; // @[Conditional.scala 39:67]
  wire  _GEN_1460 = _T_977 ? _T_1364 : spriteVisibleReg_64; // @[Conditional.scala 39:67]
  wire  _GEN_1461 = _T_977 ? _T_1365 : spriteVisibleReg_55; // @[Conditional.scala 39:67]
  wire  _GEN_1462 = _T_977 ? _T_1366 : spriteVisibleReg_63; // @[Conditional.scala 39:67]
  wire  _GEN_1463 = _T_977 ? _T_1377 : spriteVisibleReg_44; // @[Conditional.scala 39:67]
  wire  _GEN_1466 = _T_977 ? _T_1388 : spriteVisibleReg_45; // @[Conditional.scala 39:67]
  wire  _GEN_1469 = _T_977 ? _T_1399 : spriteVisibleReg_46; // @[Conditional.scala 39:67]
  wire  _GEN_1472 = _T_977 ? _T_1410 : spriteVisibleReg_47; // @[Conditional.scala 39:67]
  wire  _GEN_1475 = _T_977 ? _T_1421 : spriteVisibleReg_48; // @[Conditional.scala 39:67]
  wire  _GEN_1478 = _T_977 ? _T_1432 : spriteVisibleReg_49; // @[Conditional.scala 39:67]
  wire  _GEN_1481 = _T_977 ? _T_1443 : spriteVisibleReg_50; // @[Conditional.scala 39:67]
  wire  _GEN_1484 = _T_977 ? _T_1454 : spriteVisibleReg_51; // @[Conditional.scala 39:67]
  wire  _GEN_1488 = _T_977 ? 1'h0 : _T_1455; // @[Conditional.scala 39:67]
  wire  _GEN_1490 = _T_886 ? _GEN_1055 : spriteVisibleReg_2; // @[Conditional.scala 39:67]
  wire  _GEN_1491 = _T_886 ? _GEN_1058 : shotInteract_0; // @[Conditional.scala 39:67]
  wire  _GEN_1492 = _T_886 ? _GEN_1057 : shotPop_0; // @[Conditional.scala 39:67]
  wire  _GEN_1494 = _T_886 ? _GEN_1062 : spriteVisibleReg_3; // @[Conditional.scala 39:67]
  wire  _GEN_1495 = _T_886 ? _GEN_1064 : shotInteract_1; // @[Conditional.scala 39:67]
  wire  _GEN_1496 = _T_886 ? _GEN_1063 : shotPop_1; // @[Conditional.scala 39:67]
  wire  _GEN_1498 = _T_886 ? _GEN_1067 : spriteVisibleReg_4; // @[Conditional.scala 39:67]
  wire  _GEN_1499 = _T_886 ? _GEN_1069 : shotInteract_2; // @[Conditional.scala 39:67]
  wire  _GEN_1500 = _T_886 ? _GEN_1068 : shotPop_2; // @[Conditional.scala 39:67]
  wire  _GEN_1502 = _T_886 ? _GEN_1043 : spriteVisibleReg_5; // @[Conditional.scala 39:67]
  wire  _GEN_1503 = _T_886 ? _GEN_1046 : shotInteract_3; // @[Conditional.scala 39:67]
  wire  _GEN_1504 = _T_886 ? _GEN_1045 : shotPop_3; // @[Conditional.scala 39:67]
  wire  _GEN_1506 = _T_886 ? _GEN_1049 : spriteVisibleReg_6; // @[Conditional.scala 39:67]
  wire  _GEN_1507 = _T_886 ? _GEN_1052 : shotInteract_4; // @[Conditional.scala 39:67]
  wire  _GEN_1508 = _T_886 ? _GEN_1051 : shotPop_4; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_1517 = _T_886 ? _GEN_1059 : 2'h2; // @[Conditional.scala 39:67]
  wire  _GEN_1572 = _T_886 ? show : _GEN_1352; // @[Conditional.scala 39:67]
  wire  _GEN_1583 = _T_886 ? shipInteract : _GEN_1363; // @[Conditional.scala 39:67]
  wire  _GEN_1647 = _T_886 ? spriteVisibleReg_26 : _GEN_1427; // @[Conditional.scala 39:67]
  wire  _GEN_1650 = _T_886 ? spriteVisibleReg_30 : _GEN_1430; // @[Conditional.scala 39:67]
  wire  _GEN_1653 = _T_886 ? spriteVisibleReg_27 : _GEN_1433; // @[Conditional.scala 39:67]
  wire  _GEN_1656 = _T_886 ? spriteVisibleReg_31 : _GEN_1436; // @[Conditional.scala 39:67]
  wire  _GEN_1659 = _T_886 ? spriteVisibleReg_28 : _GEN_1439; // @[Conditional.scala 39:67]
  wire  _GEN_1662 = _T_886 ? spriteVisibleReg_32 : _GEN_1442; // @[Conditional.scala 39:67]
  wire  _GEN_1665 = _T_886 ? spriteVisibleReg_29 : _GEN_1445; // @[Conditional.scala 39:67]
  wire  _GEN_1668 = _T_886 ? spriteVisibleReg_33 : _GEN_1448; // @[Conditional.scala 39:67]
  wire  _GEN_1671 = _T_886 ? spriteVisibleReg_72 : _GEN_1451; // @[Conditional.scala 39:67]
  wire  _GEN_1672 = _T_886 ? spriteVisibleReg_66 : _GEN_1452; // @[Conditional.scala 39:67]
  wire  _GEN_1673 = _T_886 ? spriteVisibleReg_57 : _GEN_1453; // @[Conditional.scala 39:67]
  wire  _GEN_1674 = _T_886 ? spriteVisibleReg_61 : _GEN_1454; // @[Conditional.scala 39:67]
  wire  _GEN_1675 = _T_886 ? spriteVisibleReg_71 : _GEN_1455; // @[Conditional.scala 39:67]
  wire  _GEN_1676 = _T_886 ? spriteVisibleReg_65 : _GEN_1456; // @[Conditional.scala 39:67]
  wire  _GEN_1677 = _T_886 ? spriteVisibleReg_56 : _GEN_1457; // @[Conditional.scala 39:67]
  wire  _GEN_1678 = _T_886 ? spriteVisibleReg_62 : _GEN_1458; // @[Conditional.scala 39:67]
  wire  _GEN_1679 = _T_886 ? spriteVisibleReg_70 : _GEN_1459; // @[Conditional.scala 39:67]
  wire  _GEN_1680 = _T_886 ? spriteVisibleReg_64 : _GEN_1460; // @[Conditional.scala 39:67]
  wire  _GEN_1681 = _T_886 ? spriteVisibleReg_55 : _GEN_1461; // @[Conditional.scala 39:67]
  wire  _GEN_1682 = _T_886 ? spriteVisibleReg_63 : _GEN_1462; // @[Conditional.scala 39:67]
  wire  _GEN_1683 = _T_886 ? spriteVisibleReg_44 : _GEN_1463; // @[Conditional.scala 39:67]
  wire  _GEN_1686 = _T_886 ? spriteVisibleReg_45 : _GEN_1466; // @[Conditional.scala 39:67]
  wire  _GEN_1689 = _T_886 ? spriteVisibleReg_46 : _GEN_1469; // @[Conditional.scala 39:67]
  wire  _GEN_1692 = _T_886 ? spriteVisibleReg_47 : _GEN_1472; // @[Conditional.scala 39:67]
  wire  _GEN_1695 = _T_886 ? spriteVisibleReg_48 : _GEN_1475; // @[Conditional.scala 39:67]
  wire  _GEN_1698 = _T_886 ? spriteVisibleReg_49 : _GEN_1478; // @[Conditional.scala 39:67]
  wire  _GEN_1701 = _T_886 ? spriteVisibleReg_50 : _GEN_1481; // @[Conditional.scala 39:67]
  wire  _GEN_1704 = _T_886 ? spriteVisibleReg_51 : _GEN_1484; // @[Conditional.scala 39:67]
  wire  _GEN_1707 = _T_886 ? 1'h0 : _GEN_1488; // @[Conditional.scala 39:67]
  wire  _GEN_1712 = _T_862 ? spriteVisibleReg_2 : _GEN_1490; // @[Conditional.scala 39:67]
  wire  _GEN_1713 = _T_862 ? shotInteract_0 : _GEN_1491; // @[Conditional.scala 39:67]
  wire  _GEN_1714 = _T_862 ? shotPop_0 : _GEN_1492; // @[Conditional.scala 39:67]
  wire  _GEN_1716 = _T_862 ? spriteVisibleReg_3 : _GEN_1494; // @[Conditional.scala 39:67]
  wire  _GEN_1717 = _T_862 ? shotInteract_1 : _GEN_1495; // @[Conditional.scala 39:67]
  wire  _GEN_1718 = _T_862 ? shotPop_1 : _GEN_1496; // @[Conditional.scala 39:67]
  wire  _GEN_1720 = _T_862 ? spriteVisibleReg_4 : _GEN_1498; // @[Conditional.scala 39:67]
  wire  _GEN_1721 = _T_862 ? shotInteract_2 : _GEN_1499; // @[Conditional.scala 39:67]
  wire  _GEN_1722 = _T_862 ? shotPop_2 : _GEN_1500; // @[Conditional.scala 39:67]
  wire  _GEN_1724 = _T_862 ? spriteVisibleReg_5 : _GEN_1502; // @[Conditional.scala 39:67]
  wire  _GEN_1725 = _T_862 ? shotInteract_3 : _GEN_1503; // @[Conditional.scala 39:67]
  wire  _GEN_1726 = _T_862 ? shotPop_3 : _GEN_1504; // @[Conditional.scala 39:67]
  wire  _GEN_1728 = _T_862 ? spriteVisibleReg_6 : _GEN_1506; // @[Conditional.scala 39:67]
  wire  _GEN_1729 = _T_862 ? shotInteract_4 : _GEN_1507; // @[Conditional.scala 39:67]
  wire  _GEN_1730 = _T_862 ? shotPop_4 : _GEN_1508; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_1739 = _T_862 ? 2'h2 : _GEN_1517; // @[Conditional.scala 39:67]
  wire  _GEN_1793 = _T_862 ? show : _GEN_1572; // @[Conditional.scala 39:67]
  wire  _GEN_1802 = _T_862 ? shipInteract : _GEN_1583; // @[Conditional.scala 39:67]
  wire  _GEN_1866 = _T_862 ? spriteVisibleReg_26 : _GEN_1647; // @[Conditional.scala 39:67]
  wire  _GEN_1869 = _T_862 ? spriteVisibleReg_30 : _GEN_1650; // @[Conditional.scala 39:67]
  wire  _GEN_1872 = _T_862 ? spriteVisibleReg_27 : _GEN_1653; // @[Conditional.scala 39:67]
  wire  _GEN_1875 = _T_862 ? spriteVisibleReg_31 : _GEN_1656; // @[Conditional.scala 39:67]
  wire  _GEN_1878 = _T_862 ? spriteVisibleReg_28 : _GEN_1659; // @[Conditional.scala 39:67]
  wire  _GEN_1881 = _T_862 ? spriteVisibleReg_32 : _GEN_1662; // @[Conditional.scala 39:67]
  wire  _GEN_1884 = _T_862 ? spriteVisibleReg_29 : _GEN_1665; // @[Conditional.scala 39:67]
  wire  _GEN_1887 = _T_862 ? spriteVisibleReg_33 : _GEN_1668; // @[Conditional.scala 39:67]
  wire  _GEN_1890 = _T_862 ? spriteVisibleReg_72 : _GEN_1671; // @[Conditional.scala 39:67]
  wire  _GEN_1891 = _T_862 ? spriteVisibleReg_66 : _GEN_1672; // @[Conditional.scala 39:67]
  wire  _GEN_1892 = _T_862 ? spriteVisibleReg_57 : _GEN_1673; // @[Conditional.scala 39:67]
  wire  _GEN_1893 = _T_862 ? spriteVisibleReg_61 : _GEN_1674; // @[Conditional.scala 39:67]
  wire  _GEN_1894 = _T_862 ? spriteVisibleReg_71 : _GEN_1675; // @[Conditional.scala 39:67]
  wire  _GEN_1895 = _T_862 ? spriteVisibleReg_65 : _GEN_1676; // @[Conditional.scala 39:67]
  wire  _GEN_1896 = _T_862 ? spriteVisibleReg_56 : _GEN_1677; // @[Conditional.scala 39:67]
  wire  _GEN_1897 = _T_862 ? spriteVisibleReg_62 : _GEN_1678; // @[Conditional.scala 39:67]
  wire  _GEN_1898 = _T_862 ? spriteVisibleReg_70 : _GEN_1679; // @[Conditional.scala 39:67]
  wire  _GEN_1899 = _T_862 ? spriteVisibleReg_64 : _GEN_1680; // @[Conditional.scala 39:67]
  wire  _GEN_1900 = _T_862 ? spriteVisibleReg_55 : _GEN_1681; // @[Conditional.scala 39:67]
  wire  _GEN_1901 = _T_862 ? spriteVisibleReg_63 : _GEN_1682; // @[Conditional.scala 39:67]
  wire  _GEN_1902 = _T_862 ? spriteVisibleReg_44 : _GEN_1683; // @[Conditional.scala 39:67]
  wire  _GEN_1905 = _T_862 ? spriteVisibleReg_45 : _GEN_1686; // @[Conditional.scala 39:67]
  wire  _GEN_1908 = _T_862 ? spriteVisibleReg_46 : _GEN_1689; // @[Conditional.scala 39:67]
  wire  _GEN_1911 = _T_862 ? spriteVisibleReg_47 : _GEN_1692; // @[Conditional.scala 39:67]
  wire  _GEN_1914 = _T_862 ? spriteVisibleReg_48 : _GEN_1695; // @[Conditional.scala 39:67]
  wire  _GEN_1917 = _T_862 ? spriteVisibleReg_49 : _GEN_1698; // @[Conditional.scala 39:67]
  wire  _GEN_1920 = _T_862 ? spriteVisibleReg_50 : _GEN_1701; // @[Conditional.scala 39:67]
  wire  _GEN_1923 = _T_862 ? spriteVisibleReg_51 : _GEN_1704; // @[Conditional.scala 39:67]
  wire  _GEN_1926 = _T_862 ? 1'h0 : _GEN_1707; // @[Conditional.scala 39:67]
  wire  _GEN_1931 = _T_705 ? _GEN_836 : _GEN_1713; // @[Conditional.scala 39:67]
  wire  _GEN_1932 = _T_705 ? _GEN_837 : _GEN_1714; // @[Conditional.scala 39:67]
  wire  _GEN_1933 = _T_705 ? _GEN_838 : _GEN_1712; // @[Conditional.scala 39:67]
  wire  _GEN_1934 = _T_705 ? _GEN_841 : _GEN_1717; // @[Conditional.scala 39:67]
  wire  _GEN_1935 = _T_705 ? _GEN_842 : _GEN_1718; // @[Conditional.scala 39:67]
  wire  _GEN_1936 = _T_705 ? _GEN_843 : _GEN_1716; // @[Conditional.scala 39:67]
  wire  _GEN_1937 = _T_705 ? _GEN_846 : _GEN_1721; // @[Conditional.scala 39:67]
  wire  _GEN_1938 = _T_705 ? _GEN_847 : _GEN_1722; // @[Conditional.scala 39:67]
  wire  _GEN_1939 = _T_705 ? _GEN_848 : _GEN_1720; // @[Conditional.scala 39:67]
  wire  _GEN_1940 = _T_705 ? _GEN_851 : _GEN_1725; // @[Conditional.scala 39:67]
  wire  _GEN_1941 = _T_705 ? _GEN_852 : _GEN_1726; // @[Conditional.scala 39:67]
  wire  _GEN_1942 = _T_705 ? _GEN_853 : _GEN_1724; // @[Conditional.scala 39:67]
  wire  _GEN_1943 = _T_705 ? _GEN_856 : _GEN_1729; // @[Conditional.scala 39:67]
  wire  _GEN_1944 = _T_705 ? _GEN_857 : _GEN_1730; // @[Conditional.scala 39:67]
  wire  _GEN_1945 = _T_705 ? _GEN_858 : _GEN_1728; // @[Conditional.scala 39:67]
  wire  _GEN_1966 = _T_705 ? _GEN_825 : planetUp; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_1990 = _T_705 ? 2'h2 : _GEN_1739; // @[Conditional.scala 39:67]
  wire  _GEN_2030 = _T_705 ? show : _GEN_1793; // @[Conditional.scala 39:67]
  wire  _GEN_2039 = _T_705 ? shipInteract : _GEN_1802; // @[Conditional.scala 39:67]
  wire  _GEN_2102 = _T_705 ? spriteVisibleReg_26 : _GEN_1866; // @[Conditional.scala 39:67]
  wire  _GEN_2105 = _T_705 ? spriteVisibleReg_30 : _GEN_1869; // @[Conditional.scala 39:67]
  wire  _GEN_2108 = _T_705 ? spriteVisibleReg_27 : _GEN_1872; // @[Conditional.scala 39:67]
  wire  _GEN_2111 = _T_705 ? spriteVisibleReg_31 : _GEN_1875; // @[Conditional.scala 39:67]
  wire  _GEN_2114 = _T_705 ? spriteVisibleReg_28 : _GEN_1878; // @[Conditional.scala 39:67]
  wire  _GEN_2117 = _T_705 ? spriteVisibleReg_32 : _GEN_1881; // @[Conditional.scala 39:67]
  wire  _GEN_2120 = _T_705 ? spriteVisibleReg_29 : _GEN_1884; // @[Conditional.scala 39:67]
  wire  _GEN_2123 = _T_705 ? spriteVisibleReg_33 : _GEN_1887; // @[Conditional.scala 39:67]
  wire  _GEN_2126 = _T_705 ? spriteVisibleReg_72 : _GEN_1890; // @[Conditional.scala 39:67]
  wire  _GEN_2127 = _T_705 ? spriteVisibleReg_66 : _GEN_1891; // @[Conditional.scala 39:67]
  wire  _GEN_2128 = _T_705 ? spriteVisibleReg_57 : _GEN_1892; // @[Conditional.scala 39:67]
  wire  _GEN_2129 = _T_705 ? spriteVisibleReg_61 : _GEN_1893; // @[Conditional.scala 39:67]
  wire  _GEN_2130 = _T_705 ? spriteVisibleReg_71 : _GEN_1894; // @[Conditional.scala 39:67]
  wire  _GEN_2131 = _T_705 ? spriteVisibleReg_65 : _GEN_1895; // @[Conditional.scala 39:67]
  wire  _GEN_2132 = _T_705 ? spriteVisibleReg_56 : _GEN_1896; // @[Conditional.scala 39:67]
  wire  _GEN_2133 = _T_705 ? spriteVisibleReg_62 : _GEN_1897; // @[Conditional.scala 39:67]
  wire  _GEN_2134 = _T_705 ? spriteVisibleReg_70 : _GEN_1898; // @[Conditional.scala 39:67]
  wire  _GEN_2135 = _T_705 ? spriteVisibleReg_64 : _GEN_1899; // @[Conditional.scala 39:67]
  wire  _GEN_2136 = _T_705 ? spriteVisibleReg_55 : _GEN_1900; // @[Conditional.scala 39:67]
  wire  _GEN_2137 = _T_705 ? spriteVisibleReg_63 : _GEN_1901; // @[Conditional.scala 39:67]
  wire  _GEN_2138 = _T_705 ? spriteVisibleReg_44 : _GEN_1902; // @[Conditional.scala 39:67]
  wire  _GEN_2141 = _T_705 ? spriteVisibleReg_45 : _GEN_1905; // @[Conditional.scala 39:67]
  wire  _GEN_2144 = _T_705 ? spriteVisibleReg_46 : _GEN_1908; // @[Conditional.scala 39:67]
  wire  _GEN_2147 = _T_705 ? spriteVisibleReg_47 : _GEN_1911; // @[Conditional.scala 39:67]
  wire  _GEN_2150 = _T_705 ? spriteVisibleReg_48 : _GEN_1914; // @[Conditional.scala 39:67]
  wire  _GEN_2153 = _T_705 ? spriteVisibleReg_49 : _GEN_1917; // @[Conditional.scala 39:67]
  wire  _GEN_2156 = _T_705 ? spriteVisibleReg_50 : _GEN_1920; // @[Conditional.scala 39:67]
  wire  _GEN_2159 = _T_705 ? spriteVisibleReg_51 : _GEN_1923; // @[Conditional.scala 39:67]
  wire  _GEN_2162 = _T_705 ? 1'h0 : _GEN_1926; // @[Conditional.scala 39:67]
  wire  _GEN_2167 = _T_684 ? _GEN_593 : _GEN_1931; // @[Conditional.scala 39:67]
  wire  _GEN_2168 = _T_684 ? _GEN_594 : _GEN_1932; // @[Conditional.scala 39:67]
  wire  _GEN_2169 = _T_684 ? _GEN_595 : _GEN_1933; // @[Conditional.scala 39:67]
  wire  _GEN_2170 = _T_684 ? _GEN_596 : _GEN_1934; // @[Conditional.scala 39:67]
  wire  _GEN_2171 = _T_684 ? _GEN_597 : _GEN_1935; // @[Conditional.scala 39:67]
  wire  _GEN_2172 = _T_684 ? _GEN_598 : _GEN_1936; // @[Conditional.scala 39:67]
  wire  _GEN_2173 = _T_684 ? _GEN_599 : _GEN_1937; // @[Conditional.scala 39:67]
  wire  _GEN_2174 = _T_684 ? _GEN_600 : _GEN_1938; // @[Conditional.scala 39:67]
  wire  _GEN_2175 = _T_684 ? _GEN_601 : _GEN_1939; // @[Conditional.scala 39:67]
  wire  _GEN_2181 = _T_684 ? shotInteract_3 : _GEN_1940; // @[Conditional.scala 39:67]
  wire  _GEN_2182 = _T_684 ? shotPop_3 : _GEN_1941; // @[Conditional.scala 39:67]
  wire  _GEN_2183 = _T_684 ? spriteVisibleReg_5 : _GEN_1942; // @[Conditional.scala 39:67]
  wire  _GEN_2184 = _T_684 ? shotInteract_4 : _GEN_1943; // @[Conditional.scala 39:67]
  wire  _GEN_2185 = _T_684 ? shotPop_4 : _GEN_1944; // @[Conditional.scala 39:67]
  wire  _GEN_2186 = _T_684 ? spriteVisibleReg_6 : _GEN_1945; // @[Conditional.scala 39:67]
  wire  _GEN_2203 = _T_684 ? planetUp : _GEN_1966; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2226 = _T_684 ? 2'h2 : _GEN_1990; // @[Conditional.scala 39:67]
  wire  _GEN_2266 = _T_684 ? show : _GEN_2030; // @[Conditional.scala 39:67]
  wire  _GEN_2275 = _T_684 ? shipInteract : _GEN_2039; // @[Conditional.scala 39:67]
  wire  _GEN_2338 = _T_684 ? spriteVisibleReg_26 : _GEN_2102; // @[Conditional.scala 39:67]
  wire  _GEN_2341 = _T_684 ? spriteVisibleReg_30 : _GEN_2105; // @[Conditional.scala 39:67]
  wire  _GEN_2344 = _T_684 ? spriteVisibleReg_27 : _GEN_2108; // @[Conditional.scala 39:67]
  wire  _GEN_2347 = _T_684 ? spriteVisibleReg_31 : _GEN_2111; // @[Conditional.scala 39:67]
  wire  _GEN_2350 = _T_684 ? spriteVisibleReg_28 : _GEN_2114; // @[Conditional.scala 39:67]
  wire  _GEN_2353 = _T_684 ? spriteVisibleReg_32 : _GEN_2117; // @[Conditional.scala 39:67]
  wire  _GEN_2356 = _T_684 ? spriteVisibleReg_29 : _GEN_2120; // @[Conditional.scala 39:67]
  wire  _GEN_2359 = _T_684 ? spriteVisibleReg_33 : _GEN_2123; // @[Conditional.scala 39:67]
  wire  _GEN_2362 = _T_684 ? spriteVisibleReg_72 : _GEN_2126; // @[Conditional.scala 39:67]
  wire  _GEN_2363 = _T_684 ? spriteVisibleReg_66 : _GEN_2127; // @[Conditional.scala 39:67]
  wire  _GEN_2364 = _T_684 ? spriteVisibleReg_57 : _GEN_2128; // @[Conditional.scala 39:67]
  wire  _GEN_2365 = _T_684 ? spriteVisibleReg_61 : _GEN_2129; // @[Conditional.scala 39:67]
  wire  _GEN_2366 = _T_684 ? spriteVisibleReg_71 : _GEN_2130; // @[Conditional.scala 39:67]
  wire  _GEN_2367 = _T_684 ? spriteVisibleReg_65 : _GEN_2131; // @[Conditional.scala 39:67]
  wire  _GEN_2368 = _T_684 ? spriteVisibleReg_56 : _GEN_2132; // @[Conditional.scala 39:67]
  wire  _GEN_2369 = _T_684 ? spriteVisibleReg_62 : _GEN_2133; // @[Conditional.scala 39:67]
  wire  _GEN_2370 = _T_684 ? spriteVisibleReg_70 : _GEN_2134; // @[Conditional.scala 39:67]
  wire  _GEN_2371 = _T_684 ? spriteVisibleReg_64 : _GEN_2135; // @[Conditional.scala 39:67]
  wire  _GEN_2372 = _T_684 ? spriteVisibleReg_55 : _GEN_2136; // @[Conditional.scala 39:67]
  wire  _GEN_2373 = _T_684 ? spriteVisibleReg_63 : _GEN_2137; // @[Conditional.scala 39:67]
  wire  _GEN_2374 = _T_684 ? spriteVisibleReg_44 : _GEN_2138; // @[Conditional.scala 39:67]
  wire  _GEN_2377 = _T_684 ? spriteVisibleReg_45 : _GEN_2141; // @[Conditional.scala 39:67]
  wire  _GEN_2380 = _T_684 ? spriteVisibleReg_46 : _GEN_2144; // @[Conditional.scala 39:67]
  wire  _GEN_2383 = _T_684 ? spriteVisibleReg_47 : _GEN_2147; // @[Conditional.scala 39:67]
  wire  _GEN_2386 = _T_684 ? spriteVisibleReg_48 : _GEN_2150; // @[Conditional.scala 39:67]
  wire  _GEN_2389 = _T_684 ? spriteVisibleReg_49 : _GEN_2153; // @[Conditional.scala 39:67]
  wire  _GEN_2392 = _T_684 ? spriteVisibleReg_50 : _GEN_2156; // @[Conditional.scala 39:67]
  wire  _GEN_2395 = _T_684 ? spriteVisibleReg_51 : _GEN_2159; // @[Conditional.scala 39:67]
  wire  _GEN_2398 = _T_684 ? 1'h0 : _GEN_2162; // @[Conditional.scala 39:67]
  wire  _GEN_2403 = _T_627 ? _GEN_547 : _GEN_2167; // @[Conditional.scala 39:67]
  wire  _GEN_2404 = _T_627 ? _GEN_548 : _GEN_2168; // @[Conditional.scala 39:67]
  wire  _GEN_2405 = _T_627 ? _GEN_549 : _GEN_2169; // @[Conditional.scala 39:67]
  wire  _GEN_2406 = _T_627 ? _GEN_555 : _GEN_2170; // @[Conditional.scala 39:67]
  wire  _GEN_2407 = _T_627 ? _GEN_556 : _GEN_2171; // @[Conditional.scala 39:67]
  wire  _GEN_2408 = _T_627 ? _GEN_557 : _GEN_2172; // @[Conditional.scala 39:67]
  wire  _GEN_2409 = _T_627 ? _GEN_563 : _GEN_2173; // @[Conditional.scala 39:67]
  wire  _GEN_2410 = _T_627 ? _GEN_564 : _GEN_2174; // @[Conditional.scala 39:67]
  wire  _GEN_2411 = _T_627 ? _GEN_565 : _GEN_2175; // @[Conditional.scala 39:67]
  wire  _GEN_2412 = _T_627 ? _GEN_571 : _GEN_2181; // @[Conditional.scala 39:67]
  wire  _GEN_2413 = _T_627 ? _GEN_572 : _GEN_2182; // @[Conditional.scala 39:67]
  wire  _GEN_2414 = _T_627 ? _GEN_573 : _GEN_2183; // @[Conditional.scala 39:67]
  wire  _GEN_2415 = _T_627 ? _GEN_579 : _GEN_2184; // @[Conditional.scala 39:67]
  wire  _GEN_2416 = _T_627 ? _GEN_580 : _GEN_2185; // @[Conditional.scala 39:67]
  wire  _GEN_2417 = _T_627 ? _GEN_581 : _GEN_2186; // @[Conditional.scala 39:67]
  wire  _GEN_2451 = _T_627 ? planetUp : _GEN_2203; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2472 = _T_627 ? 2'h2 : _GEN_2226; // @[Conditional.scala 39:67]
  wire  _GEN_2508 = _T_627 ? show : _GEN_2266; // @[Conditional.scala 39:67]
  wire  _GEN_2517 = _T_627 ? shipInteract : _GEN_2275; // @[Conditional.scala 39:67]
  wire  _GEN_2580 = _T_627 ? spriteVisibleReg_26 : _GEN_2338; // @[Conditional.scala 39:67]
  wire  _GEN_2583 = _T_627 ? spriteVisibleReg_30 : _GEN_2341; // @[Conditional.scala 39:67]
  wire  _GEN_2586 = _T_627 ? spriteVisibleReg_27 : _GEN_2344; // @[Conditional.scala 39:67]
  wire  _GEN_2589 = _T_627 ? spriteVisibleReg_31 : _GEN_2347; // @[Conditional.scala 39:67]
  wire  _GEN_2592 = _T_627 ? spriteVisibleReg_28 : _GEN_2350; // @[Conditional.scala 39:67]
  wire  _GEN_2595 = _T_627 ? spriteVisibleReg_32 : _GEN_2353; // @[Conditional.scala 39:67]
  wire  _GEN_2598 = _T_627 ? spriteVisibleReg_29 : _GEN_2356; // @[Conditional.scala 39:67]
  wire  _GEN_2601 = _T_627 ? spriteVisibleReg_33 : _GEN_2359; // @[Conditional.scala 39:67]
  wire  _GEN_2604 = _T_627 ? spriteVisibleReg_72 : _GEN_2362; // @[Conditional.scala 39:67]
  wire  _GEN_2605 = _T_627 ? spriteVisibleReg_66 : _GEN_2363; // @[Conditional.scala 39:67]
  wire  _GEN_2606 = _T_627 ? spriteVisibleReg_57 : _GEN_2364; // @[Conditional.scala 39:67]
  wire  _GEN_2607 = _T_627 ? spriteVisibleReg_61 : _GEN_2365; // @[Conditional.scala 39:67]
  wire  _GEN_2608 = _T_627 ? spriteVisibleReg_71 : _GEN_2366; // @[Conditional.scala 39:67]
  wire  _GEN_2609 = _T_627 ? spriteVisibleReg_65 : _GEN_2367; // @[Conditional.scala 39:67]
  wire  _GEN_2610 = _T_627 ? spriteVisibleReg_56 : _GEN_2368; // @[Conditional.scala 39:67]
  wire  _GEN_2611 = _T_627 ? spriteVisibleReg_62 : _GEN_2369; // @[Conditional.scala 39:67]
  wire  _GEN_2612 = _T_627 ? spriteVisibleReg_70 : _GEN_2370; // @[Conditional.scala 39:67]
  wire  _GEN_2613 = _T_627 ? spriteVisibleReg_64 : _GEN_2371; // @[Conditional.scala 39:67]
  wire  _GEN_2614 = _T_627 ? spriteVisibleReg_55 : _GEN_2372; // @[Conditional.scala 39:67]
  wire  _GEN_2615 = _T_627 ? spriteVisibleReg_63 : _GEN_2373; // @[Conditional.scala 39:67]
  wire  _GEN_2616 = _T_627 ? spriteVisibleReg_44 : _GEN_2374; // @[Conditional.scala 39:67]
  wire  _GEN_2619 = _T_627 ? spriteVisibleReg_45 : _GEN_2377; // @[Conditional.scala 39:67]
  wire  _GEN_2622 = _T_627 ? spriteVisibleReg_46 : _GEN_2380; // @[Conditional.scala 39:67]
  wire  _GEN_2625 = _T_627 ? spriteVisibleReg_47 : _GEN_2383; // @[Conditional.scala 39:67]
  wire  _GEN_2628 = _T_627 ? spriteVisibleReg_48 : _GEN_2386; // @[Conditional.scala 39:67]
  wire  _GEN_2631 = _T_627 ? spriteVisibleReg_49 : _GEN_2389; // @[Conditional.scala 39:67]
  wire  _GEN_2634 = _T_627 ? spriteVisibleReg_50 : _GEN_2392; // @[Conditional.scala 39:67]
  wire  _GEN_2637 = _T_627 ? spriteVisibleReg_51 : _GEN_2395; // @[Conditional.scala 39:67]
  wire  _GEN_2640 = _T_627 ? 1'h0 : _GEN_2398; // @[Conditional.scala 39:67]
  wire  _GEN_2645 = _T_570 ? _GEN_397 : _GEN_2403; // @[Conditional.scala 39:67]
  wire  _GEN_2646 = _T_570 ? _GEN_398 : _GEN_2404; // @[Conditional.scala 39:67]
  wire  _GEN_2647 = _T_570 ? _GEN_399 : _GEN_2405; // @[Conditional.scala 39:67]
  wire  _GEN_2648 = _T_570 ? _GEN_405 : _GEN_2406; // @[Conditional.scala 39:67]
  wire  _GEN_2649 = _T_570 ? _GEN_406 : _GEN_2407; // @[Conditional.scala 39:67]
  wire  _GEN_2650 = _T_570 ? _GEN_407 : _GEN_2408; // @[Conditional.scala 39:67]
  wire  _GEN_2651 = _T_570 ? _GEN_413 : _GEN_2409; // @[Conditional.scala 39:67]
  wire  _GEN_2652 = _T_570 ? _GEN_414 : _GEN_2410; // @[Conditional.scala 39:67]
  wire  _GEN_2653 = _T_570 ? _GEN_415 : _GEN_2411; // @[Conditional.scala 39:67]
  wire  _GEN_2654 = _T_570 ? _GEN_421 : _GEN_2412; // @[Conditional.scala 39:67]
  wire  _GEN_2655 = _T_570 ? _GEN_422 : _GEN_2413; // @[Conditional.scala 39:67]
  wire  _GEN_2656 = _T_570 ? _GEN_423 : _GEN_2414; // @[Conditional.scala 39:67]
  wire  _GEN_2657 = _T_570 ? _GEN_429 : _GEN_2415; // @[Conditional.scala 39:67]
  wire  _GEN_2658 = _T_570 ? _GEN_430 : _GEN_2416; // @[Conditional.scala 39:67]
  wire  _GEN_2659 = _T_570 ? _GEN_431 : _GEN_2417; // @[Conditional.scala 39:67]
  wire  _GEN_2697 = _T_570 ? planetUp : _GEN_2451; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2718 = _T_570 ? 2'h2 : _GEN_2472; // @[Conditional.scala 39:67]
  wire  _GEN_2752 = _T_570 ? show : _GEN_2508; // @[Conditional.scala 39:67]
  wire  _GEN_2761 = _T_570 ? shipInteract : _GEN_2517; // @[Conditional.scala 39:67]
  wire  _GEN_2824 = _T_570 ? spriteVisibleReg_26 : _GEN_2580; // @[Conditional.scala 39:67]
  wire  _GEN_2827 = _T_570 ? spriteVisibleReg_30 : _GEN_2583; // @[Conditional.scala 39:67]
  wire  _GEN_2830 = _T_570 ? spriteVisibleReg_27 : _GEN_2586; // @[Conditional.scala 39:67]
  wire  _GEN_2833 = _T_570 ? spriteVisibleReg_31 : _GEN_2589; // @[Conditional.scala 39:67]
  wire  _GEN_2836 = _T_570 ? spriteVisibleReg_28 : _GEN_2592; // @[Conditional.scala 39:67]
  wire  _GEN_2839 = _T_570 ? spriteVisibleReg_32 : _GEN_2595; // @[Conditional.scala 39:67]
  wire  _GEN_2842 = _T_570 ? spriteVisibleReg_29 : _GEN_2598; // @[Conditional.scala 39:67]
  wire  _GEN_2845 = _T_570 ? spriteVisibleReg_33 : _GEN_2601; // @[Conditional.scala 39:67]
  wire  _GEN_2848 = _T_570 ? spriteVisibleReg_72 : _GEN_2604; // @[Conditional.scala 39:67]
  wire  _GEN_2849 = _T_570 ? spriteVisibleReg_66 : _GEN_2605; // @[Conditional.scala 39:67]
  wire  _GEN_2850 = _T_570 ? spriteVisibleReg_57 : _GEN_2606; // @[Conditional.scala 39:67]
  wire  _GEN_2851 = _T_570 ? spriteVisibleReg_61 : _GEN_2607; // @[Conditional.scala 39:67]
  wire  _GEN_2852 = _T_570 ? spriteVisibleReg_71 : _GEN_2608; // @[Conditional.scala 39:67]
  wire  _GEN_2853 = _T_570 ? spriteVisibleReg_65 : _GEN_2609; // @[Conditional.scala 39:67]
  wire  _GEN_2854 = _T_570 ? spriteVisibleReg_56 : _GEN_2610; // @[Conditional.scala 39:67]
  wire  _GEN_2855 = _T_570 ? spriteVisibleReg_62 : _GEN_2611; // @[Conditional.scala 39:67]
  wire  _GEN_2856 = _T_570 ? spriteVisibleReg_70 : _GEN_2612; // @[Conditional.scala 39:67]
  wire  _GEN_2857 = _T_570 ? spriteVisibleReg_64 : _GEN_2613; // @[Conditional.scala 39:67]
  wire  _GEN_2858 = _T_570 ? spriteVisibleReg_55 : _GEN_2614; // @[Conditional.scala 39:67]
  wire  _GEN_2859 = _T_570 ? spriteVisibleReg_63 : _GEN_2615; // @[Conditional.scala 39:67]
  wire  _GEN_2860 = _T_570 ? spriteVisibleReg_44 : _GEN_2616; // @[Conditional.scala 39:67]
  wire  _GEN_2863 = _T_570 ? spriteVisibleReg_45 : _GEN_2619; // @[Conditional.scala 39:67]
  wire  _GEN_2866 = _T_570 ? spriteVisibleReg_46 : _GEN_2622; // @[Conditional.scala 39:67]
  wire  _GEN_2869 = _T_570 ? spriteVisibleReg_47 : _GEN_2625; // @[Conditional.scala 39:67]
  wire  _GEN_2872 = _T_570 ? spriteVisibleReg_48 : _GEN_2628; // @[Conditional.scala 39:67]
  wire  _GEN_2875 = _T_570 ? spriteVisibleReg_49 : _GEN_2631; // @[Conditional.scala 39:67]
  wire  _GEN_2878 = _T_570 ? spriteVisibleReg_50 : _GEN_2634; // @[Conditional.scala 39:67]
  wire  _GEN_2881 = _T_570 ? spriteVisibleReg_51 : _GEN_2637; // @[Conditional.scala 39:67]
  wire  _GEN_2884 = _T_570 ? 1'h0 : _GEN_2640; // @[Conditional.scala 39:67]
  wire  _GEN_2889 = _T_505 ? _GEN_259 : _GEN_2645; // @[Conditional.scala 39:67]
  wire  _GEN_2890 = _T_505 ? _GEN_260 : _GEN_2646; // @[Conditional.scala 39:67]
  wire  _GEN_2891 = _T_505 ? _GEN_261 : _GEN_2647; // @[Conditional.scala 39:67]
  wire  _GEN_2892 = _T_505 ? _GEN_262 : _GEN_2648; // @[Conditional.scala 39:67]
  wire  _GEN_2893 = _T_505 ? _GEN_263 : _GEN_2649; // @[Conditional.scala 39:67]
  wire  _GEN_2894 = _T_505 ? _GEN_264 : _GEN_2650; // @[Conditional.scala 39:67]
  wire  _GEN_2895 = _T_505 ? _GEN_265 : _GEN_2651; // @[Conditional.scala 39:67]
  wire  _GEN_2896 = _T_505 ? _GEN_266 : _GEN_2652; // @[Conditional.scala 39:67]
  wire  _GEN_2897 = _T_505 ? _GEN_267 : _GEN_2653; // @[Conditional.scala 39:67]
  wire  _GEN_2898 = _T_505 ? _GEN_268 : _GEN_2654; // @[Conditional.scala 39:67]
  wire  _GEN_2899 = _T_505 ? _GEN_269 : _GEN_2655; // @[Conditional.scala 39:67]
  wire  _GEN_2900 = _T_505 ? _GEN_270 : _GEN_2656; // @[Conditional.scala 39:67]
  wire  _GEN_2901 = _T_505 ? _GEN_271 : _GEN_2657; // @[Conditional.scala 39:67]
  wire  _GEN_2902 = _T_505 ? _GEN_272 : _GEN_2658; // @[Conditional.scala 39:67]
  wire  _GEN_2903 = _T_505 ? _GEN_273 : _GEN_2659; // @[Conditional.scala 39:67]
  wire  _GEN_2941 = _T_505 ? planetUp : _GEN_2697; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2962 = _T_505 ? 2'h2 : _GEN_2718; // @[Conditional.scala 39:67]
  wire  _GEN_2996 = _T_505 ? show : _GEN_2752; // @[Conditional.scala 39:67]
  wire  _GEN_3005 = _T_505 ? shipInteract : _GEN_2761; // @[Conditional.scala 39:67]
  wire  _GEN_3068 = _T_505 ? spriteVisibleReg_26 : _GEN_2824; // @[Conditional.scala 39:67]
  wire  _GEN_3071 = _T_505 ? spriteVisibleReg_30 : _GEN_2827; // @[Conditional.scala 39:67]
  wire  _GEN_3074 = _T_505 ? spriteVisibleReg_27 : _GEN_2830; // @[Conditional.scala 39:67]
  wire  _GEN_3077 = _T_505 ? spriteVisibleReg_31 : _GEN_2833; // @[Conditional.scala 39:67]
  wire  _GEN_3080 = _T_505 ? spriteVisibleReg_28 : _GEN_2836; // @[Conditional.scala 39:67]
  wire  _GEN_3083 = _T_505 ? spriteVisibleReg_32 : _GEN_2839; // @[Conditional.scala 39:67]
  wire  _GEN_3086 = _T_505 ? spriteVisibleReg_29 : _GEN_2842; // @[Conditional.scala 39:67]
  wire  _GEN_3089 = _T_505 ? spriteVisibleReg_33 : _GEN_2845; // @[Conditional.scala 39:67]
  wire  _GEN_3092 = _T_505 ? spriteVisibleReg_72 : _GEN_2848; // @[Conditional.scala 39:67]
  wire  _GEN_3093 = _T_505 ? spriteVisibleReg_66 : _GEN_2849; // @[Conditional.scala 39:67]
  wire  _GEN_3094 = _T_505 ? spriteVisibleReg_57 : _GEN_2850; // @[Conditional.scala 39:67]
  wire  _GEN_3095 = _T_505 ? spriteVisibleReg_61 : _GEN_2851; // @[Conditional.scala 39:67]
  wire  _GEN_3096 = _T_505 ? spriteVisibleReg_71 : _GEN_2852; // @[Conditional.scala 39:67]
  wire  _GEN_3097 = _T_505 ? spriteVisibleReg_65 : _GEN_2853; // @[Conditional.scala 39:67]
  wire  _GEN_3098 = _T_505 ? spriteVisibleReg_56 : _GEN_2854; // @[Conditional.scala 39:67]
  wire  _GEN_3099 = _T_505 ? spriteVisibleReg_62 : _GEN_2855; // @[Conditional.scala 39:67]
  wire  _GEN_3100 = _T_505 ? spriteVisibleReg_70 : _GEN_2856; // @[Conditional.scala 39:67]
  wire  _GEN_3101 = _T_505 ? spriteVisibleReg_64 : _GEN_2857; // @[Conditional.scala 39:67]
  wire  _GEN_3102 = _T_505 ? spriteVisibleReg_55 : _GEN_2858; // @[Conditional.scala 39:67]
  wire  _GEN_3103 = _T_505 ? spriteVisibleReg_63 : _GEN_2859; // @[Conditional.scala 39:67]
  wire  _GEN_3104 = _T_505 ? spriteVisibleReg_44 : _GEN_2860; // @[Conditional.scala 39:67]
  wire  _GEN_3107 = _T_505 ? spriteVisibleReg_45 : _GEN_2863; // @[Conditional.scala 39:67]
  wire  _GEN_3110 = _T_505 ? spriteVisibleReg_46 : _GEN_2866; // @[Conditional.scala 39:67]
  wire  _GEN_3113 = _T_505 ? spriteVisibleReg_47 : _GEN_2869; // @[Conditional.scala 39:67]
  wire  _GEN_3116 = _T_505 ? spriteVisibleReg_48 : _GEN_2872; // @[Conditional.scala 39:67]
  wire  _GEN_3119 = _T_505 ? spriteVisibleReg_49 : _GEN_2875; // @[Conditional.scala 39:67]
  wire  _GEN_3122 = _T_505 ? spriteVisibleReg_50 : _GEN_2878; // @[Conditional.scala 39:67]
  wire  _GEN_3125 = _T_505 ? spriteVisibleReg_51 : _GEN_2881; // @[Conditional.scala 39:67]
  wire  _GEN_3128 = _T_505 ? 1'h0 : _GEN_2884; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3129 = _T_486 ? _GEN_76 : 6'h0; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3130 = _T_486 ? _GEN_101 : 13'h0; // @[Conditional.scala 39:67]
  wire  _GEN_3131 = _T_486 & _T_408; // @[Conditional.scala 39:67]
  wire  _GEN_3138 = _T_486 ? shotInteract_0 : _GEN_2889; // @[Conditional.scala 39:67]
  wire  _GEN_3139 = _T_486 ? shotPop_0 : _GEN_2890; // @[Conditional.scala 39:67]
  wire  _GEN_3140 = _T_486 ? spriteVisibleReg_2 : _GEN_2891; // @[Conditional.scala 39:67]
  wire  _GEN_3141 = _T_486 ? shotInteract_1 : _GEN_2892; // @[Conditional.scala 39:67]
  wire  _GEN_3142 = _T_486 ? shotPop_1 : _GEN_2893; // @[Conditional.scala 39:67]
  wire  _GEN_3143 = _T_486 ? spriteVisibleReg_3 : _GEN_2894; // @[Conditional.scala 39:67]
  wire  _GEN_3144 = _T_486 ? shotInteract_2 : _GEN_2895; // @[Conditional.scala 39:67]
  wire  _GEN_3145 = _T_486 ? shotPop_2 : _GEN_2896; // @[Conditional.scala 39:67]
  wire  _GEN_3146 = _T_486 ? spriteVisibleReg_4 : _GEN_2897; // @[Conditional.scala 39:67]
  wire  _GEN_3147 = _T_486 ? shotInteract_3 : _GEN_2898; // @[Conditional.scala 39:67]
  wire  _GEN_3148 = _T_486 ? shotPop_3 : _GEN_2899; // @[Conditional.scala 39:67]
  wire  _GEN_3149 = _T_486 ? spriteVisibleReg_5 : _GEN_2900; // @[Conditional.scala 39:67]
  wire  _GEN_3150 = _T_486 ? shotInteract_4 : _GEN_2901; // @[Conditional.scala 39:67]
  wire  _GEN_3151 = _T_486 ? shotPop_4 : _GEN_2902; // @[Conditional.scala 39:67]
  wire  _GEN_3152 = _T_486 ? spriteVisibleReg_6 : _GEN_2903; // @[Conditional.scala 39:67]
  wire  _GEN_3189 = _T_486 ? planetUp : _GEN_2941; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3210 = _T_486 ? 2'h2 : _GEN_2962; // @[Conditional.scala 39:67]
  wire  _GEN_3244 = _T_486 ? show : _GEN_2996; // @[Conditional.scala 39:67]
  wire  _GEN_3253 = _T_486 ? shipInteract : _GEN_3005; // @[Conditional.scala 39:67]
  wire  _GEN_3316 = _T_486 ? spriteVisibleReg_26 : _GEN_3068; // @[Conditional.scala 39:67]
  wire  _GEN_3319 = _T_486 ? spriteVisibleReg_30 : _GEN_3071; // @[Conditional.scala 39:67]
  wire  _GEN_3322 = _T_486 ? spriteVisibleReg_27 : _GEN_3074; // @[Conditional.scala 39:67]
  wire  _GEN_3325 = _T_486 ? spriteVisibleReg_31 : _GEN_3077; // @[Conditional.scala 39:67]
  wire  _GEN_3328 = _T_486 ? spriteVisibleReg_28 : _GEN_3080; // @[Conditional.scala 39:67]
  wire  _GEN_3331 = _T_486 ? spriteVisibleReg_32 : _GEN_3083; // @[Conditional.scala 39:67]
  wire  _GEN_3334 = _T_486 ? spriteVisibleReg_29 : _GEN_3086; // @[Conditional.scala 39:67]
  wire  _GEN_3337 = _T_486 ? spriteVisibleReg_33 : _GEN_3089; // @[Conditional.scala 39:67]
  wire  _GEN_3340 = _T_486 ? spriteVisibleReg_72 : _GEN_3092; // @[Conditional.scala 39:67]
  wire  _GEN_3341 = _T_486 ? spriteVisibleReg_66 : _GEN_3093; // @[Conditional.scala 39:67]
  wire  _GEN_3342 = _T_486 ? spriteVisibleReg_57 : _GEN_3094; // @[Conditional.scala 39:67]
  wire  _GEN_3343 = _T_486 ? spriteVisibleReg_61 : _GEN_3095; // @[Conditional.scala 39:67]
  wire  _GEN_3344 = _T_486 ? spriteVisibleReg_71 : _GEN_3096; // @[Conditional.scala 39:67]
  wire  _GEN_3345 = _T_486 ? spriteVisibleReg_65 : _GEN_3097; // @[Conditional.scala 39:67]
  wire  _GEN_3346 = _T_486 ? spriteVisibleReg_56 : _GEN_3098; // @[Conditional.scala 39:67]
  wire  _GEN_3347 = _T_486 ? spriteVisibleReg_62 : _GEN_3099; // @[Conditional.scala 39:67]
  wire  _GEN_3348 = _T_486 ? spriteVisibleReg_70 : _GEN_3100; // @[Conditional.scala 39:67]
  wire  _GEN_3349 = _T_486 ? spriteVisibleReg_64 : _GEN_3101; // @[Conditional.scala 39:67]
  wire  _GEN_3350 = _T_486 ? spriteVisibleReg_55 : _GEN_3102; // @[Conditional.scala 39:67]
  wire  _GEN_3351 = _T_486 ? spriteVisibleReg_63 : _GEN_3103; // @[Conditional.scala 39:67]
  wire  _GEN_3352 = _T_486 ? spriteVisibleReg_44 : _GEN_3104; // @[Conditional.scala 39:67]
  wire  _GEN_3355 = _T_486 ? spriteVisibleReg_45 : _GEN_3107; // @[Conditional.scala 39:67]
  wire  _GEN_3358 = _T_486 ? spriteVisibleReg_46 : _GEN_3110; // @[Conditional.scala 39:67]
  wire  _GEN_3361 = _T_486 ? spriteVisibleReg_47 : _GEN_3113; // @[Conditional.scala 39:67]
  wire  _GEN_3364 = _T_486 ? spriteVisibleReg_48 : _GEN_3116; // @[Conditional.scala 39:67]
  wire  _GEN_3367 = _T_486 ? spriteVisibleReg_49 : _GEN_3119; // @[Conditional.scala 39:67]
  wire  _GEN_3370 = _T_486 ? spriteVisibleReg_50 : _GEN_3122; // @[Conditional.scala 39:67]
  wire  _GEN_3373 = _T_486 ? spriteVisibleReg_51 : _GEN_3125; // @[Conditional.scala 39:67]
  wire  _GEN_3376 = _T_486 ? 1'h0 : _GEN_3128; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3380 = _T_451 ? _GEN_93 : _GEN_3129; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3381 = _T_451 ? _GEN_94 : _GEN_3130; // @[Conditional.scala 39:67]
  wire  _GEN_3382 = _T_451 ? _GEN_95 : _GEN_3131; // @[Conditional.scala 39:67]
  wire  _GEN_3388 = _T_451 ? shotInteract_0 : _GEN_3138; // @[Conditional.scala 39:67]
  wire  _GEN_3389 = _T_451 ? shotPop_0 : _GEN_3139; // @[Conditional.scala 39:67]
  wire  _GEN_3390 = _T_451 ? spriteVisibleReg_2 : _GEN_3140; // @[Conditional.scala 39:67]
  wire  _GEN_3391 = _T_451 ? shotInteract_1 : _GEN_3141; // @[Conditional.scala 39:67]
  wire  _GEN_3392 = _T_451 ? shotPop_1 : _GEN_3142; // @[Conditional.scala 39:67]
  wire  _GEN_3393 = _T_451 ? spriteVisibleReg_3 : _GEN_3143; // @[Conditional.scala 39:67]
  wire  _GEN_3394 = _T_451 ? shotInteract_2 : _GEN_3144; // @[Conditional.scala 39:67]
  wire  _GEN_3395 = _T_451 ? shotPop_2 : _GEN_3145; // @[Conditional.scala 39:67]
  wire  _GEN_3396 = _T_451 ? spriteVisibleReg_4 : _GEN_3146; // @[Conditional.scala 39:67]
  wire  _GEN_3397 = _T_451 ? shotInteract_3 : _GEN_3147; // @[Conditional.scala 39:67]
  wire  _GEN_3398 = _T_451 ? shotPop_3 : _GEN_3148; // @[Conditional.scala 39:67]
  wire  _GEN_3399 = _T_451 ? spriteVisibleReg_5 : _GEN_3149; // @[Conditional.scala 39:67]
  wire  _GEN_3400 = _T_451 ? shotInteract_4 : _GEN_3150; // @[Conditional.scala 39:67]
  wire  _GEN_3401 = _T_451 ? shotPop_4 : _GEN_3151; // @[Conditional.scala 39:67]
  wire  _GEN_3402 = _T_451 ? spriteVisibleReg_6 : _GEN_3152; // @[Conditional.scala 39:67]
  wire  _GEN_3439 = _T_451 ? planetUp : _GEN_3189; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3460 = _T_451 ? 2'h2 : _GEN_3210; // @[Conditional.scala 39:67]
  wire  _GEN_3494 = _T_451 ? show : _GEN_3244; // @[Conditional.scala 39:67]
  wire  _GEN_3503 = _T_451 ? shipInteract : _GEN_3253; // @[Conditional.scala 39:67]
  wire  _GEN_3566 = _T_451 ? spriteVisibleReg_26 : _GEN_3316; // @[Conditional.scala 39:67]
  wire  _GEN_3569 = _T_451 ? spriteVisibleReg_30 : _GEN_3319; // @[Conditional.scala 39:67]
  wire  _GEN_3572 = _T_451 ? spriteVisibleReg_27 : _GEN_3322; // @[Conditional.scala 39:67]
  wire  _GEN_3575 = _T_451 ? spriteVisibleReg_31 : _GEN_3325; // @[Conditional.scala 39:67]
  wire  _GEN_3578 = _T_451 ? spriteVisibleReg_28 : _GEN_3328; // @[Conditional.scala 39:67]
  wire  _GEN_3581 = _T_451 ? spriteVisibleReg_32 : _GEN_3331; // @[Conditional.scala 39:67]
  wire  _GEN_3584 = _T_451 ? spriteVisibleReg_29 : _GEN_3334; // @[Conditional.scala 39:67]
  wire  _GEN_3587 = _T_451 ? spriteVisibleReg_33 : _GEN_3337; // @[Conditional.scala 39:67]
  wire  _GEN_3590 = _T_451 ? spriteVisibleReg_72 : _GEN_3340; // @[Conditional.scala 39:67]
  wire  _GEN_3591 = _T_451 ? spriteVisibleReg_66 : _GEN_3341; // @[Conditional.scala 39:67]
  wire  _GEN_3592 = _T_451 ? spriteVisibleReg_57 : _GEN_3342; // @[Conditional.scala 39:67]
  wire  _GEN_3593 = _T_451 ? spriteVisibleReg_61 : _GEN_3343; // @[Conditional.scala 39:67]
  wire  _GEN_3594 = _T_451 ? spriteVisibleReg_71 : _GEN_3344; // @[Conditional.scala 39:67]
  wire  _GEN_3595 = _T_451 ? spriteVisibleReg_65 : _GEN_3345; // @[Conditional.scala 39:67]
  wire  _GEN_3596 = _T_451 ? spriteVisibleReg_56 : _GEN_3346; // @[Conditional.scala 39:67]
  wire  _GEN_3597 = _T_451 ? spriteVisibleReg_62 : _GEN_3347; // @[Conditional.scala 39:67]
  wire  _GEN_3598 = _T_451 ? spriteVisibleReg_70 : _GEN_3348; // @[Conditional.scala 39:67]
  wire  _GEN_3599 = _T_451 ? spriteVisibleReg_64 : _GEN_3349; // @[Conditional.scala 39:67]
  wire  _GEN_3600 = _T_451 ? spriteVisibleReg_55 : _GEN_3350; // @[Conditional.scala 39:67]
  wire  _GEN_3601 = _T_451 ? spriteVisibleReg_63 : _GEN_3351; // @[Conditional.scala 39:67]
  wire  _GEN_3602 = _T_451 ? spriteVisibleReg_44 : _GEN_3352; // @[Conditional.scala 39:67]
  wire  _GEN_3605 = _T_451 ? spriteVisibleReg_45 : _GEN_3355; // @[Conditional.scala 39:67]
  wire  _GEN_3608 = _T_451 ? spriteVisibleReg_46 : _GEN_3358; // @[Conditional.scala 39:67]
  wire  _GEN_3611 = _T_451 ? spriteVisibleReg_47 : _GEN_3361; // @[Conditional.scala 39:67]
  wire  _GEN_3614 = _T_451 ? spriteVisibleReg_48 : _GEN_3364; // @[Conditional.scala 39:67]
  wire  _GEN_3617 = _T_451 ? spriteVisibleReg_49 : _GEN_3367; // @[Conditional.scala 39:67]
  wire  _GEN_3620 = _T_451 ? spriteVisibleReg_50 : _GEN_3370; // @[Conditional.scala 39:67]
  wire  _GEN_3623 = _T_451 ? spriteVisibleReg_51 : _GEN_3373; // @[Conditional.scala 39:67]
  wire  _GEN_3626 = _T_451 ? 1'h0 : _GEN_3376; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3630 = _T_404 ? _GEN_67 : _GEN_3380; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3631 = _T_404 ? _GEN_68 : _GEN_3381; // @[Conditional.scala 39:67]
  wire  _GEN_3632 = _T_404 ? _GEN_69 : _GEN_3382; // @[Conditional.scala 39:67]
  wire  _GEN_3639 = _T_404 ? shotInteract_0 : _GEN_3388; // @[Conditional.scala 39:67]
  wire  _GEN_3640 = _T_404 ? shotPop_0 : _GEN_3389; // @[Conditional.scala 39:67]
  wire  _GEN_3641 = _T_404 ? spriteVisibleReg_2 : _GEN_3390; // @[Conditional.scala 39:67]
  wire  _GEN_3642 = _T_404 ? shotInteract_1 : _GEN_3391; // @[Conditional.scala 39:67]
  wire  _GEN_3643 = _T_404 ? shotPop_1 : _GEN_3392; // @[Conditional.scala 39:67]
  wire  _GEN_3644 = _T_404 ? spriteVisibleReg_3 : _GEN_3393; // @[Conditional.scala 39:67]
  wire  _GEN_3645 = _T_404 ? shotInteract_2 : _GEN_3394; // @[Conditional.scala 39:67]
  wire  _GEN_3646 = _T_404 ? shotPop_2 : _GEN_3395; // @[Conditional.scala 39:67]
  wire  _GEN_3647 = _T_404 ? spriteVisibleReg_4 : _GEN_3396; // @[Conditional.scala 39:67]
  wire  _GEN_3648 = _T_404 ? shotInteract_3 : _GEN_3397; // @[Conditional.scala 39:67]
  wire  _GEN_3649 = _T_404 ? shotPop_3 : _GEN_3398; // @[Conditional.scala 39:67]
  wire  _GEN_3650 = _T_404 ? spriteVisibleReg_5 : _GEN_3399; // @[Conditional.scala 39:67]
  wire  _GEN_3651 = _T_404 ? shotInteract_4 : _GEN_3400; // @[Conditional.scala 39:67]
  wire  _GEN_3652 = _T_404 ? shotPop_4 : _GEN_3401; // @[Conditional.scala 39:67]
  wire  _GEN_3653 = _T_404 ? spriteVisibleReg_6 : _GEN_3402; // @[Conditional.scala 39:67]
  wire  _GEN_3690 = _T_404 ? planetUp : _GEN_3439; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3711 = _T_404 ? 2'h2 : _GEN_3460; // @[Conditional.scala 39:67]
  wire  _GEN_3744 = _T_404 ? show : _GEN_3494; // @[Conditional.scala 39:67]
  wire  _GEN_3753 = _T_404 ? shipInteract : _GEN_3503; // @[Conditional.scala 39:67]
  wire  _GEN_3816 = _T_404 ? spriteVisibleReg_26 : _GEN_3566; // @[Conditional.scala 39:67]
  wire  _GEN_3819 = _T_404 ? spriteVisibleReg_30 : _GEN_3569; // @[Conditional.scala 39:67]
  wire  _GEN_3822 = _T_404 ? spriteVisibleReg_27 : _GEN_3572; // @[Conditional.scala 39:67]
  wire  _GEN_3825 = _T_404 ? spriteVisibleReg_31 : _GEN_3575; // @[Conditional.scala 39:67]
  wire  _GEN_3828 = _T_404 ? spriteVisibleReg_28 : _GEN_3578; // @[Conditional.scala 39:67]
  wire  _GEN_3831 = _T_404 ? spriteVisibleReg_32 : _GEN_3581; // @[Conditional.scala 39:67]
  wire  _GEN_3834 = _T_404 ? spriteVisibleReg_29 : _GEN_3584; // @[Conditional.scala 39:67]
  wire  _GEN_3837 = _T_404 ? spriteVisibleReg_33 : _GEN_3587; // @[Conditional.scala 39:67]
  wire  _GEN_3840 = _T_404 ? spriteVisibleReg_72 : _GEN_3590; // @[Conditional.scala 39:67]
  wire  _GEN_3841 = _T_404 ? spriteVisibleReg_66 : _GEN_3591; // @[Conditional.scala 39:67]
  wire  _GEN_3842 = _T_404 ? spriteVisibleReg_57 : _GEN_3592; // @[Conditional.scala 39:67]
  wire  _GEN_3843 = _T_404 ? spriteVisibleReg_61 : _GEN_3593; // @[Conditional.scala 39:67]
  wire  _GEN_3844 = _T_404 ? spriteVisibleReg_71 : _GEN_3594; // @[Conditional.scala 39:67]
  wire  _GEN_3845 = _T_404 ? spriteVisibleReg_65 : _GEN_3595; // @[Conditional.scala 39:67]
  wire  _GEN_3846 = _T_404 ? spriteVisibleReg_56 : _GEN_3596; // @[Conditional.scala 39:67]
  wire  _GEN_3847 = _T_404 ? spriteVisibleReg_62 : _GEN_3597; // @[Conditional.scala 39:67]
  wire  _GEN_3848 = _T_404 ? spriteVisibleReg_70 : _GEN_3598; // @[Conditional.scala 39:67]
  wire  _GEN_3849 = _T_404 ? spriteVisibleReg_64 : _GEN_3599; // @[Conditional.scala 39:67]
  wire  _GEN_3850 = _T_404 ? spriteVisibleReg_55 : _GEN_3600; // @[Conditional.scala 39:67]
  wire  _GEN_3851 = _T_404 ? spriteVisibleReg_63 : _GEN_3601; // @[Conditional.scala 39:67]
  wire  _GEN_3852 = _T_404 ? spriteVisibleReg_44 : _GEN_3602; // @[Conditional.scala 39:67]
  wire  _GEN_3855 = _T_404 ? spriteVisibleReg_45 : _GEN_3605; // @[Conditional.scala 39:67]
  wire  _GEN_3858 = _T_404 ? spriteVisibleReg_46 : _GEN_3608; // @[Conditional.scala 39:67]
  wire  _GEN_3861 = _T_404 ? spriteVisibleReg_47 : _GEN_3611; // @[Conditional.scala 39:67]
  wire  _GEN_3864 = _T_404 ? spriteVisibleReg_48 : _GEN_3614; // @[Conditional.scala 39:67]
  wire  _GEN_3867 = _T_404 ? spriteVisibleReg_49 : _GEN_3617; // @[Conditional.scala 39:67]
  wire  _GEN_3870 = _T_404 ? spriteVisibleReg_50 : _GEN_3620; // @[Conditional.scala 39:67]
  wire  _GEN_3873 = _T_404 ? spriteVisibleReg_51 : _GEN_3623; // @[Conditional.scala 39:67]
  wire  _GEN_3876 = _T_404 ? 1'h0 : _GEN_3626; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_3897 = _T_342 ? 6'h0 : _GEN_3630; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_3898 = _T_342 ? 13'h0 : _GEN_3631; // @[Conditional.scala 39:67]
  wire  _GEN_3899 = _T_342 ? 1'h0 : _GEN_3632; // @[Conditional.scala 39:67]
  wire  _GEN_3905 = _T_342 ? shotInteract_0 : _GEN_3639; // @[Conditional.scala 39:67]
  wire  _GEN_3906 = _T_342 ? shotPop_0 : _GEN_3640; // @[Conditional.scala 39:67]
  wire  _GEN_3907 = _T_342 ? spriteVisibleReg_2 : _GEN_3641; // @[Conditional.scala 39:67]
  wire  _GEN_3908 = _T_342 ? shotInteract_1 : _GEN_3642; // @[Conditional.scala 39:67]
  wire  _GEN_3909 = _T_342 ? shotPop_1 : _GEN_3643; // @[Conditional.scala 39:67]
  wire  _GEN_3910 = _T_342 ? spriteVisibleReg_3 : _GEN_3644; // @[Conditional.scala 39:67]
  wire  _GEN_3911 = _T_342 ? shotInteract_2 : _GEN_3645; // @[Conditional.scala 39:67]
  wire  _GEN_3912 = _T_342 ? shotPop_2 : _GEN_3646; // @[Conditional.scala 39:67]
  wire  _GEN_3913 = _T_342 ? spriteVisibleReg_4 : _GEN_3647; // @[Conditional.scala 39:67]
  wire  _GEN_3914 = _T_342 ? shotInteract_3 : _GEN_3648; // @[Conditional.scala 39:67]
  wire  _GEN_3915 = _T_342 ? shotPop_3 : _GEN_3649; // @[Conditional.scala 39:67]
  wire  _GEN_3916 = _T_342 ? spriteVisibleReg_5 : _GEN_3650; // @[Conditional.scala 39:67]
  wire  _GEN_3917 = _T_342 ? shotInteract_4 : _GEN_3651; // @[Conditional.scala 39:67]
  wire  _GEN_3918 = _T_342 ? shotPop_4 : _GEN_3652; // @[Conditional.scala 39:67]
  wire  _GEN_3919 = _T_342 ? spriteVisibleReg_6 : _GEN_3653; // @[Conditional.scala 39:67]
  wire  _GEN_3947 = _T_342 ? planetUp : _GEN_3690; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_3962 = _T_342 ? 2'h2 : _GEN_3711; // @[Conditional.scala 39:67]
  wire  _GEN_3995 = _T_342 ? show : _GEN_3744; // @[Conditional.scala 39:67]
  wire  _GEN_4004 = _T_342 ? shipInteract : _GEN_3753; // @[Conditional.scala 39:67]
  wire  _GEN_4067 = _T_342 ? spriteVisibleReg_26 : _GEN_3816; // @[Conditional.scala 39:67]
  wire  _GEN_4070 = _T_342 ? spriteVisibleReg_30 : _GEN_3819; // @[Conditional.scala 39:67]
  wire  _GEN_4073 = _T_342 ? spriteVisibleReg_27 : _GEN_3822; // @[Conditional.scala 39:67]
  wire  _GEN_4076 = _T_342 ? spriteVisibleReg_31 : _GEN_3825; // @[Conditional.scala 39:67]
  wire  _GEN_4079 = _T_342 ? spriteVisibleReg_28 : _GEN_3828; // @[Conditional.scala 39:67]
  wire  _GEN_4082 = _T_342 ? spriteVisibleReg_32 : _GEN_3831; // @[Conditional.scala 39:67]
  wire  _GEN_4085 = _T_342 ? spriteVisibleReg_29 : _GEN_3834; // @[Conditional.scala 39:67]
  wire  _GEN_4088 = _T_342 ? spriteVisibleReg_33 : _GEN_3837; // @[Conditional.scala 39:67]
  wire  _GEN_4091 = _T_342 ? spriteVisibleReg_72 : _GEN_3840; // @[Conditional.scala 39:67]
  wire  _GEN_4092 = _T_342 ? spriteVisibleReg_66 : _GEN_3841; // @[Conditional.scala 39:67]
  wire  _GEN_4093 = _T_342 ? spriteVisibleReg_57 : _GEN_3842; // @[Conditional.scala 39:67]
  wire  _GEN_4094 = _T_342 ? spriteVisibleReg_61 : _GEN_3843; // @[Conditional.scala 39:67]
  wire  _GEN_4095 = _T_342 ? spriteVisibleReg_71 : _GEN_3844; // @[Conditional.scala 39:67]
  wire  _GEN_4096 = _T_342 ? spriteVisibleReg_65 : _GEN_3845; // @[Conditional.scala 39:67]
  wire  _GEN_4097 = _T_342 ? spriteVisibleReg_56 : _GEN_3846; // @[Conditional.scala 39:67]
  wire  _GEN_4098 = _T_342 ? spriteVisibleReg_62 : _GEN_3847; // @[Conditional.scala 39:67]
  wire  _GEN_4099 = _T_342 ? spriteVisibleReg_70 : _GEN_3848; // @[Conditional.scala 39:67]
  wire  _GEN_4100 = _T_342 ? spriteVisibleReg_64 : _GEN_3849; // @[Conditional.scala 39:67]
  wire  _GEN_4101 = _T_342 ? spriteVisibleReg_55 : _GEN_3850; // @[Conditional.scala 39:67]
  wire  _GEN_4102 = _T_342 ? spriteVisibleReg_63 : _GEN_3851; // @[Conditional.scala 39:67]
  wire  _GEN_4103 = _T_342 ? spriteVisibleReg_44 : _GEN_3852; // @[Conditional.scala 39:67]
  wire  _GEN_4106 = _T_342 ? spriteVisibleReg_45 : _GEN_3855; // @[Conditional.scala 39:67]
  wire  _GEN_4109 = _T_342 ? spriteVisibleReg_46 : _GEN_3858; // @[Conditional.scala 39:67]
  wire  _GEN_4112 = _T_342 ? spriteVisibleReg_47 : _GEN_3861; // @[Conditional.scala 39:67]
  wire  _GEN_4115 = _T_342 ? spriteVisibleReg_48 : _GEN_3864; // @[Conditional.scala 39:67]
  wire  _GEN_4118 = _T_342 ? spriteVisibleReg_49 : _GEN_3867; // @[Conditional.scala 39:67]
  wire  _GEN_4121 = _T_342 ? spriteVisibleReg_50 : _GEN_3870; // @[Conditional.scala 39:67]
  wire  _GEN_4124 = _T_342 ? spriteVisibleReg_51 : _GEN_3873; // @[Conditional.scala 39:67]
  wire  _GEN_4127 = _T_342 ? 1'h0 : _GEN_3876; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_4148 = _T_341 ? 6'h0 : _GEN_3897; // @[Conditional.scala 40:58]
  wire [12:0] _GEN_4149 = _T_341 ? 13'h0 : _GEN_3898; // @[Conditional.scala 40:58]
  wire  _GEN_4156 = _T_341 ? shotInteract_0 : _GEN_3905; // @[Conditional.scala 40:58]
  wire  _GEN_4157 = _T_341 ? shotPop_0 : _GEN_3906; // @[Conditional.scala 40:58]
  wire  _GEN_4158 = _T_341 ? spriteVisibleReg_2 : _GEN_3907; // @[Conditional.scala 40:58]
  wire  _GEN_4159 = _T_341 ? shotInteract_1 : _GEN_3908; // @[Conditional.scala 40:58]
  wire  _GEN_4160 = _T_341 ? shotPop_1 : _GEN_3909; // @[Conditional.scala 40:58]
  wire  _GEN_4161 = _T_341 ? spriteVisibleReg_3 : _GEN_3910; // @[Conditional.scala 40:58]
  wire  _GEN_4162 = _T_341 ? shotInteract_2 : _GEN_3911; // @[Conditional.scala 40:58]
  wire  _GEN_4163 = _T_341 ? shotPop_2 : _GEN_3912; // @[Conditional.scala 40:58]
  wire  _GEN_4164 = _T_341 ? spriteVisibleReg_4 : _GEN_3913; // @[Conditional.scala 40:58]
  wire  _GEN_4165 = _T_341 ? shotInteract_3 : _GEN_3914; // @[Conditional.scala 40:58]
  wire  _GEN_4166 = _T_341 ? shotPop_3 : _GEN_3915; // @[Conditional.scala 40:58]
  wire  _GEN_4167 = _T_341 ? spriteVisibleReg_5 : _GEN_3916; // @[Conditional.scala 40:58]
  wire  _GEN_4168 = _T_341 ? shotInteract_4 : _GEN_3917; // @[Conditional.scala 40:58]
  wire  _GEN_4169 = _T_341 ? shotPop_4 : _GEN_3918; // @[Conditional.scala 40:58]
  wire  _GEN_4170 = _T_341 ? spriteVisibleReg_6 : _GEN_3919; // @[Conditional.scala 40:58]
  wire  _GEN_4198 = _T_341 ? planetUp : _GEN_3947; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_4213 = _T_341 ? 2'h2 : _GEN_3962; // @[Conditional.scala 40:58]
  wire  _GEN_4246 = _T_341 ? show : _GEN_3995; // @[Conditional.scala 40:58]
  wire  _GEN_4255 = _T_341 ? shipInteract : _GEN_4004; // @[Conditional.scala 40:58]
  wire  _GEN_4318 = _T_341 ? spriteVisibleReg_26 : _GEN_4067; // @[Conditional.scala 40:58]
  wire  _GEN_4321 = _T_341 ? spriteVisibleReg_30 : _GEN_4070; // @[Conditional.scala 40:58]
  wire  _GEN_4324 = _T_341 ? spriteVisibleReg_27 : _GEN_4073; // @[Conditional.scala 40:58]
  wire  _GEN_4327 = _T_341 ? spriteVisibleReg_31 : _GEN_4076; // @[Conditional.scala 40:58]
  wire  _GEN_4330 = _T_341 ? spriteVisibleReg_28 : _GEN_4079; // @[Conditional.scala 40:58]
  wire  _GEN_4333 = _T_341 ? spriteVisibleReg_32 : _GEN_4082; // @[Conditional.scala 40:58]
  wire  _GEN_4336 = _T_341 ? spriteVisibleReg_29 : _GEN_4085; // @[Conditional.scala 40:58]
  wire  _GEN_4339 = _T_341 ? spriteVisibleReg_33 : _GEN_4088; // @[Conditional.scala 40:58]
  wire  _GEN_4342 = _T_341 ? spriteVisibleReg_72 : _GEN_4091; // @[Conditional.scala 40:58]
  wire  _GEN_4343 = _T_341 ? spriteVisibleReg_66 : _GEN_4092; // @[Conditional.scala 40:58]
  wire  _GEN_4344 = _T_341 ? spriteVisibleReg_57 : _GEN_4093; // @[Conditional.scala 40:58]
  wire  _GEN_4345 = _T_341 ? spriteVisibleReg_61 : _GEN_4094; // @[Conditional.scala 40:58]
  wire  _GEN_4346 = _T_341 ? spriteVisibleReg_71 : _GEN_4095; // @[Conditional.scala 40:58]
  wire  _GEN_4347 = _T_341 ? spriteVisibleReg_65 : _GEN_4096; // @[Conditional.scala 40:58]
  wire  _GEN_4348 = _T_341 ? spriteVisibleReg_56 : _GEN_4097; // @[Conditional.scala 40:58]
  wire  _GEN_4349 = _T_341 ? spriteVisibleReg_62 : _GEN_4098; // @[Conditional.scala 40:58]
  wire  _GEN_4350 = _T_341 ? spriteVisibleReg_70 : _GEN_4099; // @[Conditional.scala 40:58]
  wire  _GEN_4351 = _T_341 ? spriteVisibleReg_64 : _GEN_4100; // @[Conditional.scala 40:58]
  wire  _GEN_4352 = _T_341 ? spriteVisibleReg_55 : _GEN_4101; // @[Conditional.scala 40:58]
  wire  _GEN_4353 = _T_341 ? spriteVisibleReg_63 : _GEN_4102; // @[Conditional.scala 40:58]
  wire  _GEN_4354 = _T_341 ? spriteVisibleReg_44 : _GEN_4103; // @[Conditional.scala 40:58]
  wire  _GEN_4357 = _T_341 ? spriteVisibleReg_45 : _GEN_4106; // @[Conditional.scala 40:58]
  wire  _GEN_4360 = _T_341 ? spriteVisibleReg_46 : _GEN_4109; // @[Conditional.scala 40:58]
  wire  _GEN_4363 = _T_341 ? spriteVisibleReg_47 : _GEN_4112; // @[Conditional.scala 40:58]
  wire  _GEN_4366 = _T_341 ? spriteVisibleReg_48 : _GEN_4115; // @[Conditional.scala 40:58]
  wire  _GEN_4369 = _T_341 ? spriteVisibleReg_49 : _GEN_4118; // @[Conditional.scala 40:58]
  wire  _GEN_4372 = _T_341 ? spriteVisibleReg_50 : _GEN_4121; // @[Conditional.scala 40:58]
  wire  _GEN_4375 = _T_341 ? spriteVisibleReg_51 : _GEN_4124; // @[Conditional.scala 40:58]
  BoxDetection boxDetection ( // @[GameLogic.scala 700:28]
    .clock(boxDetection_clock),
    .io_boxXPosition_0(boxDetection_io_boxXPosition_0),
    .io_boxXPosition_2(boxDetection_io_boxXPosition_2),
    .io_boxXPosition_3(boxDetection_io_boxXPosition_3),
    .io_boxXPosition_4(boxDetection_io_boxXPosition_4),
    .io_boxXPosition_5(boxDetection_io_boxXPosition_5),
    .io_boxXPosition_6(boxDetection_io_boxXPosition_6),
    .io_boxXPosition_7(boxDetection_io_boxXPosition_7),
    .io_boxXPosition_8(boxDetection_io_boxXPosition_8),
    .io_boxXPosition_9(boxDetection_io_boxXPosition_9),
    .io_boxXPosition_10(boxDetection_io_boxXPosition_10),
    .io_boxXPosition_11(boxDetection_io_boxXPosition_11),
    .io_boxXPosition_12(boxDetection_io_boxXPosition_12),
    .io_boxXPosition_13(boxDetection_io_boxXPosition_13),
    .io_boxXPosition_14(boxDetection_io_boxXPosition_14),
    .io_boxXPosition_15(boxDetection_io_boxXPosition_15),
    .io_boxXPosition_16(boxDetection_io_boxXPosition_16),
    .io_boxXPosition_17(boxDetection_io_boxXPosition_17),
    .io_boxYPosition_0(boxDetection_io_boxYPosition_0),
    .io_boxYPosition_2(boxDetection_io_boxYPosition_2),
    .io_boxYPosition_3(boxDetection_io_boxYPosition_3),
    .io_boxYPosition_4(boxDetection_io_boxYPosition_4),
    .io_boxYPosition_5(boxDetection_io_boxYPosition_5),
    .io_boxYPosition_6(boxDetection_io_boxYPosition_6),
    .io_boxYPosition_7(boxDetection_io_boxYPosition_7),
    .io_boxYPosition_8(boxDetection_io_boxYPosition_8),
    .io_boxYPosition_9(boxDetection_io_boxYPosition_9),
    .io_boxYPosition_10(boxDetection_io_boxYPosition_10),
    .io_boxYPosition_11(boxDetection_io_boxYPosition_11),
    .io_boxYPosition_12(boxDetection_io_boxYPosition_12),
    .io_boxYPosition_13(boxDetection_io_boxYPosition_13),
    .io_boxYPosition_14(boxDetection_io_boxYPosition_14),
    .io_boxYPosition_15(boxDetection_io_boxYPosition_15),
    .io_boxYPosition_16(boxDetection_io_boxYPosition_16),
    .io_boxYPosition_17(boxDetection_io_boxYPosition_17),
    .io_overlap_0_7(boxDetection_io_overlap_0_7),
    .io_overlap_0_8(boxDetection_io_overlap_0_8),
    .io_overlap_0_9(boxDetection_io_overlap_0_9),
    .io_overlap_0_10(boxDetection_io_overlap_0_10),
    .io_overlap_0_11(boxDetection_io_overlap_0_11),
    .io_overlap_0_12(boxDetection_io_overlap_0_12),
    .io_overlap_0_13(boxDetection_io_overlap_0_13),
    .io_overlap_0_14(boxDetection_io_overlap_0_14),
    .io_overlap_0_15(boxDetection_io_overlap_0_15),
    .io_overlap_0_16(boxDetection_io_overlap_0_16),
    .io_overlap_0_17(boxDetection_io_overlap_0_17),
    .io_overlap_2_7(boxDetection_io_overlap_2_7),
    .io_overlap_2_8(boxDetection_io_overlap_2_8),
    .io_overlap_2_9(boxDetection_io_overlap_2_9),
    .io_overlap_2_10(boxDetection_io_overlap_2_10),
    .io_overlap_2_11(boxDetection_io_overlap_2_11),
    .io_overlap_2_12(boxDetection_io_overlap_2_12),
    .io_overlap_2_13(boxDetection_io_overlap_2_13),
    .io_overlap_2_14(boxDetection_io_overlap_2_14),
    .io_overlap_2_15(boxDetection_io_overlap_2_15),
    .io_overlap_2_16(boxDetection_io_overlap_2_16),
    .io_overlap_2_17(boxDetection_io_overlap_2_17),
    .io_overlap_3_7(boxDetection_io_overlap_3_7),
    .io_overlap_3_8(boxDetection_io_overlap_3_8),
    .io_overlap_3_9(boxDetection_io_overlap_3_9),
    .io_overlap_3_10(boxDetection_io_overlap_3_10),
    .io_overlap_3_11(boxDetection_io_overlap_3_11),
    .io_overlap_3_12(boxDetection_io_overlap_3_12),
    .io_overlap_3_13(boxDetection_io_overlap_3_13),
    .io_overlap_3_14(boxDetection_io_overlap_3_14),
    .io_overlap_3_15(boxDetection_io_overlap_3_15),
    .io_overlap_3_16(boxDetection_io_overlap_3_16),
    .io_overlap_3_17(boxDetection_io_overlap_3_17),
    .io_overlap_4_7(boxDetection_io_overlap_4_7),
    .io_overlap_4_8(boxDetection_io_overlap_4_8),
    .io_overlap_4_9(boxDetection_io_overlap_4_9),
    .io_overlap_4_10(boxDetection_io_overlap_4_10),
    .io_overlap_4_11(boxDetection_io_overlap_4_11),
    .io_overlap_4_12(boxDetection_io_overlap_4_12),
    .io_overlap_4_13(boxDetection_io_overlap_4_13),
    .io_overlap_4_14(boxDetection_io_overlap_4_14),
    .io_overlap_4_15(boxDetection_io_overlap_4_15),
    .io_overlap_4_16(boxDetection_io_overlap_4_16),
    .io_overlap_4_17(boxDetection_io_overlap_4_17),
    .io_overlap_5_7(boxDetection_io_overlap_5_7),
    .io_overlap_5_8(boxDetection_io_overlap_5_8),
    .io_overlap_5_9(boxDetection_io_overlap_5_9),
    .io_overlap_5_10(boxDetection_io_overlap_5_10),
    .io_overlap_5_11(boxDetection_io_overlap_5_11),
    .io_overlap_5_12(boxDetection_io_overlap_5_12),
    .io_overlap_5_13(boxDetection_io_overlap_5_13),
    .io_overlap_5_14(boxDetection_io_overlap_5_14),
    .io_overlap_5_15(boxDetection_io_overlap_5_15),
    .io_overlap_5_16(boxDetection_io_overlap_5_16),
    .io_overlap_5_17(boxDetection_io_overlap_5_17),
    .io_overlap_6_7(boxDetection_io_overlap_6_7),
    .io_overlap_6_8(boxDetection_io_overlap_6_8),
    .io_overlap_6_9(boxDetection_io_overlap_6_9),
    .io_overlap_6_10(boxDetection_io_overlap_6_10),
    .io_overlap_6_11(boxDetection_io_overlap_6_11),
    .io_overlap_6_12(boxDetection_io_overlap_6_12),
    .io_overlap_6_13(boxDetection_io_overlap_6_13),
    .io_overlap_6_14(boxDetection_io_overlap_6_14),
    .io_overlap_6_15(boxDetection_io_overlap_6_15),
    .io_overlap_6_17(boxDetection_io_overlap_6_17)
  );
  Randomizer Randomizer ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_clock),
    .reset(Randomizer_reset),
    .io_out(Randomizer_io_out)
  );
  Randomizer_1 Randomizer_1 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_1_clock),
    .reset(Randomizer_1_reset),
    .io_out(Randomizer_1_io_out)
  );
  Randomizer_2 Randomizer_2 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_2_clock),
    .reset(Randomizer_2_reset),
    .io_out(Randomizer_2_io_out)
  );
  Randomizer_3 Randomizer_3 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_3_clock),
    .reset(Randomizer_3_reset),
    .io_out(Randomizer_3_io_out)
  );
  Randomizer_4 Randomizer_4 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_4_clock),
    .reset(Randomizer_4_reset),
    .io_out(Randomizer_4_io_out)
  );
  Randomizer_5 Randomizer_5 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_5_clock),
    .reset(Randomizer_5_reset),
    .io_out(Randomizer_5_io_out)
  );
  Randomizer_6 Randomizer_6 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_6_clock),
    .reset(Randomizer_6_reset),
    .io_out(Randomizer_6_io_out)
  );
  Randomizer_7 Randomizer_7 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_7_clock),
    .reset(Randomizer_7_reset),
    .io_out(Randomizer_7_io_out)
  );
  Randomizer_8 Randomizer_8 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_8_clock),
    .reset(Randomizer_8_reset),
    .io_out(Randomizer_8_io_out)
  );
  Randomizer_9 Randomizer_9 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_9_clock),
    .reset(Randomizer_9_reset),
    .io_out(Randomizer_9_io_out)
  );
  Randomizer_10 Randomizer_10 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_10_clock),
    .reset(Randomizer_10_reset),
    .io_out(Randomizer_10_io_out)
  );
  Randomizer_11 Randomizer_11 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_11_clock),
    .reset(Randomizer_11_reset),
    .io_out(Randomizer_11_io_out)
  );
  Randomizer_12 Randomizer_12 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_12_clock),
    .reset(Randomizer_12_reset),
    .io_out(Randomizer_12_io_out)
  );
  Randomizer_13 Randomizer_13 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_13_clock),
    .reset(Randomizer_13_reset),
    .io_out(Randomizer_13_io_out)
  );
  Randomizer_14 Randomizer_14 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_14_clock),
    .reset(Randomizer_14_reset),
    .io_out(Randomizer_14_io_out)
  );
  Randomizer_15 Randomizer_15 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_15_clock),
    .reset(Randomizer_15_reset),
    .io_out(Randomizer_15_io_out)
  );
  Randomizer_16 Randomizer_16 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_16_clock),
    .reset(Randomizer_16_reset),
    .io_out(Randomizer_16_io_out)
  );
  Randomizer_17 Randomizer_17 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_17_clock),
    .reset(Randomizer_17_reset),
    .io_out(Randomizer_17_io_out)
  );
  Randomizer_18 Randomizer_18 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_18_clock),
    .reset(Randomizer_18_reset),
    .io_out(Randomizer_18_io_out)
  );
  Randomizer_19 Randomizer_19 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_19_clock),
    .reset(Randomizer_19_reset),
    .io_out(Randomizer_19_io_out)
  );
  Randomizer Randomizer_20 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_20_clock),
    .reset(Randomizer_20_reset),
    .io_out(Randomizer_20_io_out)
  );
  Randomizer_1 Randomizer_21 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_21_clock),
    .reset(Randomizer_21_reset),
    .io_out(Randomizer_21_io_out)
  );
  Randomizer_2 Randomizer_22 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_22_clock),
    .reset(Randomizer_22_reset),
    .io_out(Randomizer_22_io_out)
  );
  Randomizer_3 Randomizer_23 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_23_clock),
    .reset(Randomizer_23_reset),
    .io_out(Randomizer_23_io_out)
  );
  Randomizer_4 Randomizer_24 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_24_clock),
    .reset(Randomizer_24_reset),
    .io_out(Randomizer_24_io_out)
  );
  Randomizer_5 Randomizer_25 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_25_clock),
    .reset(Randomizer_25_reset),
    .io_out(Randomizer_25_io_out)
  );
  Randomizer_8 Randomizer_26 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_26_clock),
    .reset(Randomizer_26_reset),
    .io_out(Randomizer_26_io_out)
  );
  Randomizer_9 Randomizer_27 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_27_clock),
    .reset(Randomizer_27_reset),
    .io_out(Randomizer_27_io_out)
  );
  Randomizer_10 Randomizer_28 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_28_clock),
    .reset(Randomizer_28_reset),
    .io_out(Randomizer_28_io_out)
  );
  Randomizer_11 Randomizer_29 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_29_clock),
    .reset(Randomizer_29_reset),
    .io_out(Randomizer_29_io_out)
  );
  Randomizer_18 Randomizer_30 ( // @[GameLogic.scala 189:24]
    .clock(Randomizer_30_clock),
    .reset(Randomizer_30_reset),
    .io_out(Randomizer_30_io_out)
  );
  Randomizer_19 Randomizer_31 ( // @[GameLogic.scala 190:31]
    .clock(Randomizer_31_clock),
    .reset(Randomizer_31_reset),
    .io_out(Randomizer_31_io_out)
  );
  Randomizer_4 Randomizer_32 ( // @[GameLogic.scala 362:24]
    .clock(Randomizer_32_clock),
    .reset(Randomizer_32_reset),
    .io_out(Randomizer_32_io_out)
  );
  Randomizer_33 Randomizer_33 ( // @[GameLogic.scala 118:24]
    .clock(Randomizer_33_clock),
    .reset(Randomizer_33_reset),
    .io_out(Randomizer_33_io_out)
  );
  Randomizer_34 Randomizer_34 ( // @[GameLogic.scala 95:24]
    .clock(Randomizer_34_clock),
    .reset(Randomizer_34_reset),
    .io_out(Randomizer_34_io_out)
  );
  Randomizer_35 Randomizer_35 ( // @[GameLogic.scala 96:25]
    .clock(Randomizer_35_clock),
    .reset(Randomizer_35_reset),
    .io_out(Randomizer_35_io_out)
  );
  Randomizer_36 Randomizer_36 ( // @[GameLogic.scala 95:24]
    .clock(Randomizer_36_clock),
    .reset(Randomizer_36_reset),
    .io_out(Randomizer_36_io_out)
  );
  Randomizer_35 Randomizer_37 ( // @[GameLogic.scala 96:25]
    .clock(Randomizer_37_clock),
    .reset(Randomizer_37_reset),
    .io_out(Randomizer_37_io_out)
  );
  Randomizer_38 Randomizer_38 ( // @[GameLogic.scala 95:24]
    .clock(Randomizer_38_clock),
    .reset(Randomizer_38_reset),
    .io_out(Randomizer_38_io_out)
  );
  Randomizer_35 Randomizer_39 ( // @[GameLogic.scala 96:25]
    .clock(Randomizer_39_clock),
    .reset(Randomizer_39_reset),
    .io_out(Randomizer_39_io_out)
  );
  Randomizer_40 Randomizer_40 ( // @[GameLogic.scala 118:24]
    .clock(Randomizer_40_clock),
    .reset(Randomizer_40_reset),
    .io_out(Randomizer_40_io_out)
  );
  Randomizer_41 Randomizer_41 ( // @[GameLogic.scala 95:24]
    .clock(Randomizer_41_clock),
    .reset(Randomizer_41_reset),
    .io_out(Randomizer_41_io_out)
  );
  Randomizer_35 Randomizer_42 ( // @[GameLogic.scala 96:25]
    .clock(Randomizer_42_clock),
    .reset(Randomizer_42_reset),
    .io_out(Randomizer_42_io_out)
  );
  Randomizer_43 Randomizer_43 ( // @[GameLogic.scala 95:24]
    .clock(Randomizer_43_clock),
    .reset(Randomizer_43_reset),
    .io_out(Randomizer_43_io_out)
  );
  Randomizer_35 Randomizer_44 ( // @[GameLogic.scala 96:25]
    .clock(Randomizer_44_clock),
    .reset(Randomizer_44_reset),
    .io_out(Randomizer_44_io_out)
  );
  Randomizer_45 Randomizer_45 ( // @[GameLogic.scala 95:24]
    .clock(Randomizer_45_clock),
    .reset(Randomizer_45_reset),
    .io_out(Randomizer_45_io_out)
  );
  Randomizer_35 Randomizer_46 ( // @[GameLogic.scala 96:25]
    .clock(Randomizer_46_clock),
    .reset(Randomizer_46_reset),
    .io_out(Randomizer_46_io_out)
  );
  assign io_songInput = {{2'd0}, _GEN_4213}; // @[GameLogic.scala 51:16 GameLogic.scala 221:21 GameLogic.scala 221:21 GameLogic.scala 221:21]
  assign io_spriteXPosition_0 = Xstart_0; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_1 = Xstart_1; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_2 = Xstart_2; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_3 = Xstart_3; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_4 = Xstart_4; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_5 = Xstart_5; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_6 = Xstart_6; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_7 = Xstart_7; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_8 = Xstart_8; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_9 = Xstart_9; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_10 = Xstart_10; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_11 = Xstart_11; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_12 = Xstart_12; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_13 = Xstart_13; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_14 = Xstart_14; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_15 = Xstart_15; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_16 = Xstart_16; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_17 = Xstart_17; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_18 = Xstart_18; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_19 = Xstart_19; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_20 = Xstart_20; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_21 = Xstart_21; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_22 = Xstart_22; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_23 = Xstart_23; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_24 = Xstart_24; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_25 = Xstart_25; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_26 = Xstart_26; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_27 = Xstart_27; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_28 = Xstart_28; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_29 = Xstart_29; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_30 = Xstart_30; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_31 = Xstart_31; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_32 = Xstart_32; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_33 = Xstart_33; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_41 = Xstart_41; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_42 = Xstart_42; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_43 = Xstart_43; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_44 = Xstart_44; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_45 = Xstart_45; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_46 = Xstart_46; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_47 = Xstart_47; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_48 = Xstart_48; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_49 = Xstart_49; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_50 = Xstart_50; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_51 = Xstart_51; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_122 = Xstart_122; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_123 = Xstart_123; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_124 = Xstart_124; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_125 = Xstart_125; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_126 = Xstart_126; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteXPosition_127 = Xstart_127; // @[GameLogic.scala 57:22 GameLogic.scala 627:27]
  assign io_spriteYPosition_0 = Ystart_0[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_1 = Ystart_1[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_2 = Ystart_2[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_3 = Ystart_3[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_4 = Ystart_4[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_5 = Ystart_5[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_6 = Ystart_6[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_7 = Ystart_7[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_8 = Ystart_8[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_9 = Ystart_9[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_10 = Ystart_10[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_11 = Ystart_11[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_12 = Ystart_12[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_13 = Ystart_13[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_14 = Ystart_14[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_15 = Ystart_15[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_16 = Ystart_16[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_17 = Ystart_17[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_18 = Ystart_18[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_19 = Ystart_19[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_20 = Ystart_20[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_21 = Ystart_21[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_22 = Ystart_22[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_23 = Ystart_23[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_24 = Ystart_24[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_25 = Ystart_25[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_26 = Ystart_26[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_27 = Ystart_27[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_28 = Ystart_28[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_29 = Ystart_29[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_30 = Ystart_30[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_31 = Ystart_31[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_32 = Ystart_32[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_33 = Ystart_33[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_41 = Ystart_41[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_42 = Ystart_42[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_43 = Ystart_43[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_122 = Ystart_122[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_123 = Ystart_123[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_124 = Ystart_124[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_125 = Ystart_125[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_126 = Ystart_126[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteYPosition_127 = Ystart_127[9:0]; // @[GameLogic.scala 58:22 GameLogic.scala 628:27]
  assign io_spriteVisible_0 = _T_281 ? 1'h0 : spriteVisibleReg_0; // @[GameLogic.scala 59:20 GameLogic.scala 629:25 GameLogic.scala 331:27]
  assign io_spriteVisible_1 = _T_281 ? 1'h0 : spriteVisibleReg_1; // @[GameLogic.scala 59:20 GameLogic.scala 629:25 GameLogic.scala 332:27]
  assign io_spriteVisible_2 = spriteVisibleReg_2; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_3 = spriteVisibleReg_3; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_4 = spriteVisibleReg_4; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_5 = spriteVisibleReg_5; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_6 = spriteVisibleReg_6; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_7 = spriteVisibleReg_7; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_8 = spriteVisibleReg_8; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_9 = spriteVisibleReg_9; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_10 = spriteVisibleReg_10; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_11 = spriteVisibleReg_11; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_12 = spriteVisibleReg_12; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_13 = spriteVisibleReg_13; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_14 = spriteVisibleReg_14; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_15 = spriteVisibleReg_15; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_16 = spriteVisibleReg_16; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_17 = spriteVisibleReg_17; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_18 = spriteVisibleReg_18; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_19 = spriteVisibleReg_19; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_20 = spriteVisibleReg_20; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_21 = spriteVisibleReg_21; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_22 = spriteVisibleReg_22; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_23 = spriteVisibleReg_23; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_24 = spriteVisibleReg_24; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_25 = spriteVisibleReg_25; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_26 = spriteVisibleReg_26; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_27 = spriteVisibleReg_27; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_28 = spriteVisibleReg_28; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_29 = spriteVisibleReg_29; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_30 = spriteVisibleReg_30; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_31 = spriteVisibleReg_31; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_32 = spriteVisibleReg_32; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_33 = spriteVisibleReg_33; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_41 = spriteVisibleReg_41; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_42 = spriteVisibleReg_42; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_43 = spriteVisibleReg_43; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_44 = spriteVisibleReg_44; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_45 = spriteVisibleReg_45; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_46 = spriteVisibleReg_46; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_47 = spriteVisibleReg_47; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_48 = spriteVisibleReg_48; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_49 = spriteVisibleReg_49; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_50 = spriteVisibleReg_50; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_51 = spriteVisibleReg_51; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_55 = spriteVisibleReg_55; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_56 = spriteVisibleReg_56; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_57 = spriteVisibleReg_57; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_61 = spriteVisibleReg_61; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_62 = spriteVisibleReg_62; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_63 = spriteVisibleReg_63; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_64 = spriteVisibleReg_64; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_65 = spriteVisibleReg_65; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_66 = spriteVisibleReg_66; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_70 = spriteVisibleReg_70; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_71 = spriteVisibleReg_71; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteVisible_72 = spriteVisibleReg_72; // @[GameLogic.scala 59:20 GameLogic.scala 629:25]
  assign io_spriteFlipVertical_122 = spriteFlipVerticalReg_122; // @[GameLogic.scala 61:25 GameLogic.scala 631:30]
  assign io_spriteFlipVertical_123 = spriteFlipVerticalReg_123; // @[GameLogic.scala 61:25 GameLogic.scala 631:30]
  assign io_spriteFlipVertical_124 = spriteFlipVerticalReg_124; // @[GameLogic.scala 61:25 GameLogic.scala 631:30]
  assign io_spriteFlipVertical_125 = spriteFlipVerticalReg_125; // @[GameLogic.scala 61:25 GameLogic.scala 631:30]
  assign io_spriteFlipVertical_126 = spriteFlipVerticalReg_126; // @[GameLogic.scala 61:25 GameLogic.scala 631:30]
  assign io_spriteFlipVertical_127 = spriteFlipVerticalReg_127; // @[GameLogic.scala 61:25 GameLogic.scala 631:30]
  assign io_viewBoxX_0 = viewX; // @[GameLogic.scala 633:15 GameLogic.scala 638:18]
  assign io_backBufferWriteData = _GEN_4148[4:0]; // @[GameLogic.scala 642:26 GameLogic.scala 757:36 GameLogic.scala 773:34 GameLogic.scala 787:34 GameLogic.scala 809:34 GameLogic.scala 822:34 GameLogic.scala 836:32]
  assign io_backBufferWriteAddress = _GEN_4149[10:0]; // @[GameLogic.scala 643:29 GameLogic.scala 758:39 GameLogic.scala 774:37 GameLogic.scala 788:37 GameLogic.scala 810:37 GameLogic.scala 823:37 GameLogic.scala 837:35]
  assign io_backBufferWriteEnable = _T_341 ? 1'h0 : _GEN_3899; // @[GameLogic.scala 644:28 GameLogic.scala 759:38 GameLogic.scala 775:36 GameLogic.scala 789:36 GameLogic.scala 811:36 GameLogic.scala 824:36 GameLogic.scala 838:34]
  assign io_frameUpdateDone = _T_341 ? 1'h0 : _GEN_4127; // @[GameLogic.scala 647:22 GameLogic.scala 1025:26]
  assign boxDetection_clock = clock;
  assign boxDetection_io_boxXPosition_0 = $signed(Xstart_0) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_2 = $signed(Xstart_2) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_3 = $signed(Xstart_3) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_4 = $signed(Xstart_4) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_5 = $signed(Xstart_5) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_6 = $signed(Xstart_6) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_7 = $signed(Xstart_7) + $signed(_GEN_4393); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_8 = $signed(Xstart_8) + $signed(_GEN_4395); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_9 = $signed(Xstart_9) + $signed(_GEN_4397); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_10 = $signed(Xstart_10) + $signed(_GEN_4397); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_11 = $signed(Xstart_11) + $signed(_GEN_4397); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_12 = $signed(Xstart_12) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_13 = $signed(Xstart_13) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_14 = $signed(Xstart_14) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_15 = $signed(Xstart_15) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_16 = $signed(Xstart_16) + $signed(_GEN_4379); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxXPosition_17 = $signed(Xstart_17) + $signed(_GEN_4413); // @[GameLogic.scala 702:35]
  assign boxDetection_io_boxYPosition_0 = _T_42[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_2 = _T_70[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_3 = _T_84[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_4 = _T_98[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_5 = _T_112[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_6 = _T_126[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_7 = _T_140[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_8 = _T_154[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_9 = _T_168[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_10 = _T_182[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_11 = _T_196[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_12 = _T_210[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_13 = _T_224[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_14 = _T_238[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_15 = _T_252[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_16 = _T_266[9:0]; // @[GameLogic.scala 703:35]
  assign boxDetection_io_boxYPosition_17 = _T_280[9:0]; // @[GameLogic.scala 703:35]
  assign Randomizer_clock = clock;
  assign Randomizer_reset = reset;
  assign Randomizer_1_clock = clock;
  assign Randomizer_1_reset = reset;
  assign Randomizer_2_clock = clock;
  assign Randomizer_2_reset = reset;
  assign Randomizer_3_clock = clock;
  assign Randomizer_3_reset = reset;
  assign Randomizer_4_clock = clock;
  assign Randomizer_4_reset = reset;
  assign Randomizer_5_clock = clock;
  assign Randomizer_5_reset = reset;
  assign Randomizer_6_clock = clock;
  assign Randomizer_6_reset = reset;
  assign Randomizer_7_clock = clock;
  assign Randomizer_7_reset = reset;
  assign Randomizer_8_clock = clock;
  assign Randomizer_8_reset = reset;
  assign Randomizer_9_clock = clock;
  assign Randomizer_9_reset = reset;
  assign Randomizer_10_clock = clock;
  assign Randomizer_10_reset = reset;
  assign Randomizer_11_clock = clock;
  assign Randomizer_11_reset = reset;
  assign Randomizer_12_clock = clock;
  assign Randomizer_12_reset = reset;
  assign Randomizer_13_clock = clock;
  assign Randomizer_13_reset = reset;
  assign Randomizer_14_clock = clock;
  assign Randomizer_14_reset = reset;
  assign Randomizer_15_clock = clock;
  assign Randomizer_15_reset = reset;
  assign Randomizer_16_clock = clock;
  assign Randomizer_16_reset = reset;
  assign Randomizer_17_clock = clock;
  assign Randomizer_17_reset = reset;
  assign Randomizer_18_clock = clock;
  assign Randomizer_18_reset = reset;
  assign Randomizer_19_clock = clock;
  assign Randomizer_19_reset = reset;
  assign Randomizer_20_clock = clock;
  assign Randomizer_20_reset = reset;
  assign Randomizer_21_clock = clock;
  assign Randomizer_21_reset = reset;
  assign Randomizer_22_clock = clock;
  assign Randomizer_22_reset = reset;
  assign Randomizer_23_clock = clock;
  assign Randomizer_23_reset = reset;
  assign Randomizer_24_clock = clock;
  assign Randomizer_24_reset = reset;
  assign Randomizer_25_clock = clock;
  assign Randomizer_25_reset = reset;
  assign Randomizer_26_clock = clock;
  assign Randomizer_26_reset = reset;
  assign Randomizer_27_clock = clock;
  assign Randomizer_27_reset = reset;
  assign Randomizer_28_clock = clock;
  assign Randomizer_28_reset = reset;
  assign Randomizer_29_clock = clock;
  assign Randomizer_29_reset = reset;
  assign Randomizer_30_clock = clock;
  assign Randomizer_30_reset = reset;
  assign Randomizer_31_clock = clock;
  assign Randomizer_31_reset = reset;
  assign Randomizer_32_clock = clock;
  assign Randomizer_32_reset = reset;
  assign Randomizer_33_clock = clock;
  assign Randomizer_33_reset = reset;
  assign Randomizer_34_clock = clock;
  assign Randomizer_34_reset = reset;
  assign Randomizer_35_clock = clock;
  assign Randomizer_35_reset = reset;
  assign Randomizer_36_clock = clock;
  assign Randomizer_36_reset = reset;
  assign Randomizer_37_clock = clock;
  assign Randomizer_37_reset = reset;
  assign Randomizer_38_clock = clock;
  assign Randomizer_38_reset = reset;
  assign Randomizer_39_clock = clock;
  assign Randomizer_39_reset = reset;
  assign Randomizer_40_clock = clock;
  assign Randomizer_40_reset = reset;
  assign Randomizer_41_clock = clock;
  assign Randomizer_41_reset = reset;
  assign Randomizer_42_clock = clock;
  assign Randomizer_42_reset = reset;
  assign Randomizer_43_clock = clock;
  assign Randomizer_43_reset = reset;
  assign Randomizer_44_clock = clock;
  assign Randomizer_44_reset = reset;
  assign Randomizer_45_clock = clock;
  assign Randomizer_45_reset = reset;
  assign Randomizer_46_clock = clock;
  assign Randomizer_46_reset = reset;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  planetUp = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  Xstart_0 = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  Xstart_1 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  Xstart_2 = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  Xstart_3 = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  Xstart_4 = _RAND_5[10:0];
  _RAND_6 = {1{`RANDOM}};
  Xstart_5 = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  Xstart_6 = _RAND_7[10:0];
  _RAND_8 = {1{`RANDOM}};
  Xstart_7 = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  Xstart_8 = _RAND_9[10:0];
  _RAND_10 = {1{`RANDOM}};
  Xstart_9 = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  Xstart_10 = _RAND_11[10:0];
  _RAND_12 = {1{`RANDOM}};
  Xstart_11 = _RAND_12[10:0];
  _RAND_13 = {1{`RANDOM}};
  Xstart_12 = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  Xstart_13 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  Xstart_14 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  Xstart_15 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  Xstart_16 = _RAND_17[10:0];
  _RAND_18 = {1{`RANDOM}};
  Xstart_17 = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  Xstart_18 = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  Xstart_19 = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  Xstart_20 = _RAND_21[10:0];
  _RAND_22 = {1{`RANDOM}};
  Xstart_21 = _RAND_22[10:0];
  _RAND_23 = {1{`RANDOM}};
  Xstart_22 = _RAND_23[10:0];
  _RAND_24 = {1{`RANDOM}};
  Xstart_23 = _RAND_24[10:0];
  _RAND_25 = {1{`RANDOM}};
  Xstart_24 = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  Xstart_25 = _RAND_26[10:0];
  _RAND_27 = {1{`RANDOM}};
  Xstart_26 = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  Xstart_27 = _RAND_28[10:0];
  _RAND_29 = {1{`RANDOM}};
  Xstart_28 = _RAND_29[10:0];
  _RAND_30 = {1{`RANDOM}};
  Xstart_29 = _RAND_30[10:0];
  _RAND_31 = {1{`RANDOM}};
  Xstart_30 = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  Xstart_31 = _RAND_32[10:0];
  _RAND_33 = {1{`RANDOM}};
  Xstart_32 = _RAND_33[10:0];
  _RAND_34 = {1{`RANDOM}};
  Xstart_33 = _RAND_34[10:0];
  _RAND_35 = {1{`RANDOM}};
  Xstart_41 = _RAND_35[10:0];
  _RAND_36 = {1{`RANDOM}};
  Xstart_42 = _RAND_36[10:0];
  _RAND_37 = {1{`RANDOM}};
  Xstart_43 = _RAND_37[10:0];
  _RAND_38 = {1{`RANDOM}};
  Xstart_44 = _RAND_38[10:0];
  _RAND_39 = {1{`RANDOM}};
  Xstart_45 = _RAND_39[10:0];
  _RAND_40 = {1{`RANDOM}};
  Xstart_46 = _RAND_40[10:0];
  _RAND_41 = {1{`RANDOM}};
  Xstart_47 = _RAND_41[10:0];
  _RAND_42 = {1{`RANDOM}};
  Xstart_48 = _RAND_42[10:0];
  _RAND_43 = {1{`RANDOM}};
  Xstart_49 = _RAND_43[10:0];
  _RAND_44 = {1{`RANDOM}};
  Xstart_50 = _RAND_44[10:0];
  _RAND_45 = {1{`RANDOM}};
  Xstart_51 = _RAND_45[10:0];
  _RAND_46 = {1{`RANDOM}};
  Xstart_122 = _RAND_46[10:0];
  _RAND_47 = {1{`RANDOM}};
  Xstart_123 = _RAND_47[10:0];
  _RAND_48 = {1{`RANDOM}};
  Xstart_124 = _RAND_48[10:0];
  _RAND_49 = {1{`RANDOM}};
  Xstart_125 = _RAND_49[10:0];
  _RAND_50 = {1{`RANDOM}};
  Xstart_126 = _RAND_50[10:0];
  _RAND_51 = {1{`RANDOM}};
  Xstart_127 = _RAND_51[10:0];
  _RAND_52 = {1{`RANDOM}};
  Ystart_0 = _RAND_52[10:0];
  _RAND_53 = {1{`RANDOM}};
  Ystart_1 = _RAND_53[10:0];
  _RAND_54 = {1{`RANDOM}};
  Ystart_2 = _RAND_54[10:0];
  _RAND_55 = {1{`RANDOM}};
  Ystart_3 = _RAND_55[10:0];
  _RAND_56 = {1{`RANDOM}};
  Ystart_4 = _RAND_56[10:0];
  _RAND_57 = {1{`RANDOM}};
  Ystart_5 = _RAND_57[10:0];
  _RAND_58 = {1{`RANDOM}};
  Ystart_6 = _RAND_58[10:0];
  _RAND_59 = {1{`RANDOM}};
  Ystart_7 = _RAND_59[10:0];
  _RAND_60 = {1{`RANDOM}};
  Ystart_8 = _RAND_60[10:0];
  _RAND_61 = {1{`RANDOM}};
  Ystart_9 = _RAND_61[10:0];
  _RAND_62 = {1{`RANDOM}};
  Ystart_10 = _RAND_62[10:0];
  _RAND_63 = {1{`RANDOM}};
  Ystart_11 = _RAND_63[10:0];
  _RAND_64 = {1{`RANDOM}};
  Ystart_12 = _RAND_64[10:0];
  _RAND_65 = {1{`RANDOM}};
  Ystart_13 = _RAND_65[10:0];
  _RAND_66 = {1{`RANDOM}};
  Ystart_14 = _RAND_66[10:0];
  _RAND_67 = {1{`RANDOM}};
  Ystart_15 = _RAND_67[10:0];
  _RAND_68 = {1{`RANDOM}};
  Ystart_16 = _RAND_68[10:0];
  _RAND_69 = {1{`RANDOM}};
  Ystart_17 = _RAND_69[10:0];
  _RAND_70 = {1{`RANDOM}};
  Ystart_18 = _RAND_70[10:0];
  _RAND_71 = {1{`RANDOM}};
  Ystart_19 = _RAND_71[10:0];
  _RAND_72 = {1{`RANDOM}};
  Ystart_20 = _RAND_72[10:0];
  _RAND_73 = {1{`RANDOM}};
  Ystart_21 = _RAND_73[10:0];
  _RAND_74 = {1{`RANDOM}};
  Ystart_22 = _RAND_74[10:0];
  _RAND_75 = {1{`RANDOM}};
  Ystart_23 = _RAND_75[10:0];
  _RAND_76 = {1{`RANDOM}};
  Ystart_24 = _RAND_76[10:0];
  _RAND_77 = {1{`RANDOM}};
  Ystart_25 = _RAND_77[10:0];
  _RAND_78 = {1{`RANDOM}};
  Ystart_26 = _RAND_78[10:0];
  _RAND_79 = {1{`RANDOM}};
  Ystart_27 = _RAND_79[10:0];
  _RAND_80 = {1{`RANDOM}};
  Ystart_28 = _RAND_80[10:0];
  _RAND_81 = {1{`RANDOM}};
  Ystart_29 = _RAND_81[10:0];
  _RAND_82 = {1{`RANDOM}};
  Ystart_30 = _RAND_82[10:0];
  _RAND_83 = {1{`RANDOM}};
  Ystart_31 = _RAND_83[10:0];
  _RAND_84 = {1{`RANDOM}};
  Ystart_32 = _RAND_84[10:0];
  _RAND_85 = {1{`RANDOM}};
  Ystart_33 = _RAND_85[10:0];
  _RAND_86 = {1{`RANDOM}};
  Ystart_41 = _RAND_86[10:0];
  _RAND_87 = {1{`RANDOM}};
  Ystart_42 = _RAND_87[10:0];
  _RAND_88 = {1{`RANDOM}};
  Ystart_43 = _RAND_88[10:0];
  _RAND_89 = {1{`RANDOM}};
  Ystart_122 = _RAND_89[10:0];
  _RAND_90 = {1{`RANDOM}};
  Ystart_123 = _RAND_90[10:0];
  _RAND_91 = {1{`RANDOM}};
  Ystart_124 = _RAND_91[10:0];
  _RAND_92 = {1{`RANDOM}};
  Ystart_125 = _RAND_92[10:0];
  _RAND_93 = {1{`RANDOM}};
  Ystart_126 = _RAND_93[10:0];
  _RAND_94 = {1{`RANDOM}};
  Ystart_127 = _RAND_94[10:0];
  _RAND_95 = {1{`RANDOM}};
  spriteVisibleReg_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  spriteVisibleReg_1 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  spriteVisibleReg_2 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  spriteVisibleReg_3 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  spriteVisibleReg_4 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  spriteVisibleReg_5 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  spriteVisibleReg_6 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  spriteVisibleReg_7 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  spriteVisibleReg_8 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  spriteVisibleReg_9 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  spriteVisibleReg_10 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  spriteVisibleReg_11 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  spriteVisibleReg_12 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  spriteVisibleReg_13 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  spriteVisibleReg_14 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  spriteVisibleReg_15 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  spriteVisibleReg_16 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  spriteVisibleReg_17 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  spriteVisibleReg_18 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  spriteVisibleReg_19 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  spriteVisibleReg_20 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  spriteVisibleReg_21 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  spriteVisibleReg_22 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  spriteVisibleReg_23 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  spriteVisibleReg_24 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  spriteVisibleReg_25 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  spriteVisibleReg_26 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  spriteVisibleReg_27 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  spriteVisibleReg_28 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  spriteVisibleReg_29 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  spriteVisibleReg_30 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  spriteVisibleReg_31 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  spriteVisibleReg_32 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  spriteVisibleReg_33 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  spriteVisibleReg_41 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  spriteVisibleReg_42 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  spriteVisibleReg_43 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  spriteVisibleReg_44 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  spriteVisibleReg_45 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  spriteVisibleReg_46 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  spriteVisibleReg_47 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  spriteVisibleReg_48 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  spriteVisibleReg_49 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  spriteVisibleReg_50 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  spriteVisibleReg_51 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  spriteVisibleReg_55 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  spriteVisibleReg_56 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  spriteVisibleReg_57 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  spriteVisibleReg_61 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  spriteVisibleReg_62 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  spriteVisibleReg_63 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  spriteVisibleReg_64 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  spriteVisibleReg_65 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  spriteVisibleReg_66 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  spriteVisibleReg_70 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  spriteVisibleReg_71 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  spriteVisibleReg_72 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  spriteFlipVerticalReg_122 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  spriteFlipVerticalReg_123 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  spriteFlipVerticalReg_124 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  spriteFlipVerticalReg_125 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  spriteFlipVerticalReg_126 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  spriteFlipVerticalReg_127 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  btnCReg = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  viewX = _RAND_159[9:0];
  _RAND_160 = {1{`RANDOM}};
  stateReg = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  shotCnt = _RAND_161[9:0];
  _RAND_162 = {1{`RANDOM}};
  shotLoad = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  shotCntBig = _RAND_163[2:0];
  _RAND_164 = {1{`RANDOM}};
  shotCntFast = _RAND_164[2:0];
  _RAND_165 = {1{`RANDOM}};
  shotPop_0 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  shotPop_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  shotPop_2 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  shotPop_3 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  shotPop_4 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  shotInteract_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  shotInteract_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  shotInteract_2 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  shotInteract_3 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  shotInteract_4 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  astInteract_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  astInteract_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  astInteract_2 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  astInteract_3 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  astInteract_4 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  astInteract_5 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  astInteract_6 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  astInteract_7 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  astInteract_8 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  astInteract_9 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  astInteract_10 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  shipInteract = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  die_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  die_1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  die_2 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  die_3 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  die_4 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  die_5 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  die_6 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  die_7 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  die_8 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  die_9 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  die_10 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  kill_0_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  kill_0_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  kill_0_2 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  kill_0_3 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  kill_0_4 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  kill_1_0 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  kill_1_1 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  kill_1_2 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  kill_1_3 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  kill_1_4 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  kill_2_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  kill_2_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  kill_2_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  kill_2_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  kill_2_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  kill_3_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  kill_3_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  kill_3_2 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  kill_3_3 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  kill_3_4 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  kill_4_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  kill_4_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  kill_4_2 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  kill_4_3 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  kill_4_4 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  kill_5_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  kill_5_1 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  kill_5_2 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  kill_5_3 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  kill_5_4 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  kill_6_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  kill_6_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  kill_6_2 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  kill_6_3 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  kill_6_4 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  kill_7_0 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  kill_7_1 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  kill_7_2 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  kill_7_3 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  kill_7_4 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  kill_8_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  kill_8_1 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  kill_8_2 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  kill_8_3 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  kill_8_4 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  kill_9_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  kill_9_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  kill_9_2 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  kill_9_3 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  kill_10_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  kill_10_1 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  kill_10_2 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  kill_10_3 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  kill_10_4 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  hp = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  planetHp = _RAND_253[4:0];
  _RAND_254 = {1{`RANDOM}};
  spwnProt = _RAND_254[5:0];
  _RAND_255 = {1{`RANDOM}};
  show = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  blink = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  secCnt = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  level = _RAND_258[2:0];
  _RAND_259 = {1{`RANDOM}};
  start = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  levelCng = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  cngCnt = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  cnt = _RAND_262[9:0];
  _RAND_263 = {1{`RANDOM}};
  count1 = _RAND_263[6:0];
  _RAND_264 = {1{`RANDOM}};
  count3 = _RAND_264[6:0];
  _RAND_265 = {1{`RANDOM}};
  count4 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  count5 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  _T_912 = _RAND_267[10:0];
  _RAND_268 = {1{`RANDOM}};
  _T_917 = _RAND_268[10:0];
  _RAND_269 = {1{`RANDOM}};
  _T_927 = _RAND_269[10:0];
  _RAND_270 = {1{`RANDOM}};
  _T_932 = _RAND_270[10:0];
  _RAND_271 = {1{`RANDOM}};
  _T_940 = _RAND_271[10:0];
  _RAND_272 = {1{`RANDOM}};
  _T_945 = _RAND_272[10:0];
  _RAND_273 = {1{`RANDOM}};
  _T_953 = _RAND_273[10:0];
  _RAND_274 = {1{`RANDOM}};
  _T_958 = _RAND_274[10:0];
  _RAND_275 = {1{`RANDOM}};
  _T_966 = _RAND_275[10:0];
  _RAND_276 = {1{`RANDOM}};
  _T_971 = _RAND_276[10:0];
  _RAND_277 = {1{`RANDOM}};
  _T_978 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_979 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  _T_980 = _RAND_279[2:0];
  _RAND_280 = {1{`RANDOM}};
  _T_981 = _RAND_280[2:0];
  _RAND_281 = {1{`RANDOM}};
  _T_982 = _RAND_281[2:0];
  _RAND_282 = {1{`RANDOM}};
  _T_1028 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  _T_1029 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_1030 = _RAND_284[2:0];
  _RAND_285 = {1{`RANDOM}};
  _T_1031 = _RAND_285[2:0];
  _RAND_286 = {1{`RANDOM}};
  _T_1032 = _RAND_286[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    planetUp <= reset | _GEN_4198;
    if (reset) begin
      Xstart_0 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (_T_862) begin
                          if (_T_863) begin
                            if (io_btnR) begin
                              if (_T_875) begin
                                Xstart_0 <= _T_878;
                              end
                            end else if (io_btnL) begin
                              if (_T_882) begin
                                Xstart_0 <= _T_885;
                              end
                            end
                          end
                        end else if (!(_T_886)) begin
                          if (_T_977) begin
                            if (die_10) begin
                              if (_T_1134) begin
                                Xstart_0 <= 11'sh40;
                              end else if (die_9) begin
                                if (_T_1134) begin
                                  Xstart_0 <= 11'sh40;
                                end else if (die_8) begin
                                  if (_T_1134) begin
                                    Xstart_0 <= 11'sh40;
                                  end else if (die_7) begin
                                    if (_T_1134) begin
                                      Xstart_0 <= 11'sh40;
                                    end else if (die_6) begin
                                      if (_T_1134) begin
                                        Xstart_0 <= 11'sh40;
                                      end else if (die_5) begin
                                        if (_T_1134) begin
                                          Xstart_0 <= 11'sh40;
                                        end else if (die_4) begin
                                          if (_T_1134) begin
                                            Xstart_0 <= 11'sh40;
                                          end else if (die_3) begin
                                            if (_T_1134) begin
                                              Xstart_0 <= 11'sh40;
                                            end else if (die_2) begin
                                              if (_T_1134) begin
                                                Xstart_0 <= 11'sh40;
                                              end else if (die_1) begin
                                                if (_T_1134) begin
                                                  Xstart_0 <= 11'sh40;
                                                end else if (die_0) begin
                                                  if (_T_1134) begin
                                                    Xstart_0 <= 11'sh40;
                                                  end
                                                end
                                              end else if (die_0) begin
                                                if (_T_1134) begin
                                                  Xstart_0 <= 11'sh40;
                                                end
                                              end
                                            end else if (die_1) begin
                                              if (_T_1134) begin
                                                Xstart_0 <= 11'sh40;
                                              end else if (die_0) begin
                                                if (_T_1134) begin
                                                  Xstart_0 <= 11'sh40;
                                                end
                                              end
                                            end else if (die_0) begin
                                              if (_T_1134) begin
                                                Xstart_0 <= 11'sh40;
                                              end
                                            end
                                          end else if (die_2) begin
                                            if (_T_1134) begin
                                              Xstart_0 <= 11'sh40;
                                            end else if (die_1) begin
                                              if (_T_1134) begin
                                                Xstart_0 <= 11'sh40;
                                              end else begin
                                                Xstart_0 <= _GEN_1182;
                                              end
                                            end else begin
                                              Xstart_0 <= _GEN_1182;
                                            end
                                          end else if (die_1) begin
                                            if (_T_1134) begin
                                              Xstart_0 <= 11'sh40;
                                            end else begin
                                              Xstart_0 <= _GEN_1182;
                                            end
                                          end else begin
                                            Xstart_0 <= _GEN_1182;
                                          end
                                        end else if (die_3) begin
                                          if (_T_1134) begin
                                            Xstart_0 <= 11'sh40;
                                          end else if (die_2) begin
                                            if (_T_1134) begin
                                              Xstart_0 <= 11'sh40;
                                            end else begin
                                              Xstart_0 <= _GEN_1192;
                                            end
                                          end else begin
                                            Xstart_0 <= _GEN_1192;
                                          end
                                        end else if (die_2) begin
                                          if (_T_1134) begin
                                            Xstart_0 <= 11'sh40;
                                          end else begin
                                            Xstart_0 <= _GEN_1192;
                                          end
                                        end else begin
                                          Xstart_0 <= _GEN_1192;
                                        end
                                      end else if (die_4) begin
                                        if (_T_1134) begin
                                          Xstart_0 <= 11'sh40;
                                        end else if (die_3) begin
                                          if (_T_1134) begin
                                            Xstart_0 <= 11'sh40;
                                          end else begin
                                            Xstart_0 <= _GEN_1202;
                                          end
                                        end else begin
                                          Xstart_0 <= _GEN_1202;
                                        end
                                      end else if (die_3) begin
                                        if (_T_1134) begin
                                          Xstart_0 <= 11'sh40;
                                        end else begin
                                          Xstart_0 <= _GEN_1202;
                                        end
                                      end else begin
                                        Xstart_0 <= _GEN_1202;
                                      end
                                    end else if (die_5) begin
                                      if (_T_1134) begin
                                        Xstart_0 <= 11'sh40;
                                      end else if (die_4) begin
                                        if (_T_1134) begin
                                          Xstart_0 <= 11'sh40;
                                        end else begin
                                          Xstart_0 <= _GEN_1212;
                                        end
                                      end else begin
                                        Xstart_0 <= _GEN_1212;
                                      end
                                    end else if (die_4) begin
                                      if (_T_1134) begin
                                        Xstart_0 <= 11'sh40;
                                      end else begin
                                        Xstart_0 <= _GEN_1212;
                                      end
                                    end else begin
                                      Xstart_0 <= _GEN_1212;
                                    end
                                  end else if (die_6) begin
                                    if (_T_1134) begin
                                      Xstart_0 <= 11'sh40;
                                    end else if (die_5) begin
                                      if (_T_1134) begin
                                        Xstart_0 <= 11'sh40;
                                      end else begin
                                        Xstart_0 <= _GEN_1222;
                                      end
                                    end else begin
                                      Xstart_0 <= _GEN_1222;
                                    end
                                  end else if (die_5) begin
                                    if (_T_1134) begin
                                      Xstart_0 <= 11'sh40;
                                    end else begin
                                      Xstart_0 <= _GEN_1222;
                                    end
                                  end else begin
                                    Xstart_0 <= _GEN_1222;
                                  end
                                end else if (die_7) begin
                                  if (_T_1134) begin
                                    Xstart_0 <= 11'sh40;
                                  end else if (die_6) begin
                                    if (_T_1134) begin
                                      Xstart_0 <= 11'sh40;
                                    end else begin
                                      Xstart_0 <= _GEN_1232;
                                    end
                                  end else begin
                                    Xstart_0 <= _GEN_1232;
                                  end
                                end else if (die_6) begin
                                  if (_T_1134) begin
                                    Xstart_0 <= 11'sh40;
                                  end else begin
                                    Xstart_0 <= _GEN_1232;
                                  end
                                end else begin
                                  Xstart_0 <= _GEN_1232;
                                end
                              end else if (die_8) begin
                                if (_T_1134) begin
                                  Xstart_0 <= 11'sh40;
                                end else if (die_7) begin
                                  if (_T_1134) begin
                                    Xstart_0 <= 11'sh40;
                                  end else begin
                                    Xstart_0 <= _GEN_1242;
                                  end
                                end else begin
                                  Xstart_0 <= _GEN_1242;
                                end
                              end else if (die_7) begin
                                if (_T_1134) begin
                                  Xstart_0 <= 11'sh40;
                                end else begin
                                  Xstart_0 <= _GEN_1242;
                                end
                              end else begin
                                Xstart_0 <= _GEN_1242;
                              end
                            end else if (die_9) begin
                              if (_T_1134) begin
                                Xstart_0 <= 11'sh40;
                              end else if (die_8) begin
                                if (_T_1134) begin
                                  Xstart_0 <= 11'sh40;
                                end else begin
                                  Xstart_0 <= _GEN_1252;
                                end
                              end else begin
                                Xstart_0 <= _GEN_1252;
                              end
                            end else if (die_8) begin
                              if (_T_1134) begin
                                Xstart_0 <= 11'sh40;
                              end else begin
                                Xstart_0 <= _GEN_1252;
                              end
                            end else begin
                              Xstart_0 <= _GEN_1252;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_1 <= 11'sh20;
    end else begin
      Xstart_1 <= Xstart_0;
    end
    if (reset) begin
      Xstart_2 <= 11'sh258;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_2 <= _T_348;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (!(_T_705)) begin
                      if (!(_T_862)) begin
                        if (_T_886) begin
                          if (_T_863) begin
                            if (_T_909) begin
                              Xstart_2 <= _T_889;
                            end else if (_T_924) begin
                              Xstart_2 <= _T_889;
                            end else if (shotPop_0) begin
                              if (shotLoad) begin
                                Xstart_2 <= _T_944;
                              end else begin
                                Xstart_2 <= _T_889;
                              end
                            end else begin
                              Xstart_2 <= _T_889;
                            end
                          end else begin
                            Xstart_2 <= _T_889;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_3 <= 11'sh258;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_3 <= _T_351;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (!(_T_705)) begin
                      if (!(_T_862)) begin
                        if (_T_886) begin
                          if (_T_863) begin
                            if (_T_909) begin
                              Xstart_3 <= _T_893;
                            end else if (_T_924) begin
                              Xstart_3 <= _T_893;
                            end else if (shotPop_0) begin
                              Xstart_3 <= _T_893;
                            end else if (shotPop_1) begin
                              if (shotLoad) begin
                                Xstart_3 <= _T_957;
                              end else begin
                                Xstart_3 <= _T_893;
                              end
                            end else begin
                              Xstart_3 <= _T_893;
                            end
                          end else begin
                            Xstart_3 <= _T_893;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_4 <= 11'sh258;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_4 <= _T_354;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (!(_T_705)) begin
                      if (!(_T_862)) begin
                        if (_T_886) begin
                          if (_T_863) begin
                            if (_T_909) begin
                              Xstart_4 <= _T_897;
                            end else if (_T_924) begin
                              Xstart_4 <= _T_897;
                            end else if (shotPop_0) begin
                              Xstart_4 <= _T_897;
                            end else if (shotPop_1) begin
                              Xstart_4 <= _T_897;
                            end else if (shotPop_2) begin
                              if (shotLoad) begin
                                Xstart_4 <= _T_970;
                              end else begin
                                Xstart_4 <= _T_897;
                              end
                            end else begin
                              Xstart_4 <= _T_897;
                            end
                          end else begin
                            Xstart_4 <= _T_897;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_5 <= 11'sh258;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_5 <= _T_357;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (!(_T_705)) begin
                      if (!(_T_862)) begin
                        if (_T_886) begin
                          if (_T_863) begin
                            if (_T_909) begin
                              if (shotPop_3) begin
                                if (shotLoad) begin
                                  Xstart_5 <= _T_916;
                                end else begin
                                  Xstart_5 <= _T_901;
                                end
                              end else begin
                                Xstart_5 <= _T_901;
                              end
                            end else begin
                              Xstart_5 <= _T_901;
                            end
                          end else begin
                            Xstart_5 <= _T_901;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_6 <= 11'sh258;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_6 <= _T_360;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (!(_T_705)) begin
                      if (!(_T_862)) begin
                        if (_T_886) begin
                          if (_T_863) begin
                            if (_T_909) begin
                              Xstart_6 <= _T_905;
                            end else if (_T_924) begin
                              if (shotPop_4) begin
                                if (shotLoad) begin
                                  Xstart_6 <= _T_931;
                                end else begin
                                  Xstart_6 <= _T_905;
                                end
                              end else begin
                                Xstart_6 <= _T_905;
                              end
                            end else begin
                              Xstart_6 <= _T_905;
                            end
                          end else begin
                            Xstart_6 <= _T_905;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_7 <= 11'sh226;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_7 <= _T_363;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (_T_505) begin
              if (_T_507) begin
                if (_T_511) begin
                  if (_T_514) begin
                    if (_T_501) begin
                      Xstart_7 <= _T_294;
                    end else begin
                      Xstart_7 <= _T_525;
                    end
                  end else begin
                    Xstart_7 <= _T_510;
                  end
                end else begin
                  Xstart_7 <= _T_510;
                end
              end
            end else if (!(_T_570)) begin
              if (!(_T_627)) begin
                if (!(_T_684)) begin
                  if (_T_705) begin
                    if (_T_706) begin
                      if (_T_511) begin
                        if (_T_514) begin
                          if (_T_501) begin
                            Xstart_7 <= _T_294;
                          end else begin
                            Xstart_7 <= _T_525;
                          end
                        end else begin
                          Xstart_7 <= _T_510;
                        end
                      end else begin
                        Xstart_7 <= _T_510;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_8 <= 11'sh262;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_8 <= _T_366;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (_T_505) begin
              if (_T_507) begin
                if (_T_511) begin
                  if (_T_532) begin
                    if (_T_501) begin
                      Xstart_8 <= _T_294;
                    end else begin
                      Xstart_8 <= _T_525;
                    end
                  end else begin
                    Xstart_8 <= _T_528;
                  end
                end else begin
                  Xstart_8 <= _T_528;
                end
              end
            end else if (!(_T_570)) begin
              if (!(_T_627)) begin
                if (!(_T_684)) begin
                  if (_T_705) begin
                    if (_T_706) begin
                      if (_T_511) begin
                        if (_T_532) begin
                          if (_T_501) begin
                            Xstart_8 <= _T_294;
                          end else begin
                            Xstart_8 <= _T_525;
                          end
                        end else begin
                          Xstart_8 <= _T_528;
                        end
                      end else begin
                        Xstart_8 <= _T_528;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_9 <= 11'sh320;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_9 <= _T_369;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (_T_505) begin
              if (_T_507) begin
                if (_T_511) begin
                  if (_T_550) begin
                    Xstart_9 <= _GEN_105;
                  end else begin
                    Xstart_9 <= _T_546;
                  end
                end else begin
                  Xstart_9 <= _T_546;
                end
              end
            end else if (!(_T_570)) begin
              if (!(_T_627)) begin
                if (!(_T_684)) begin
                  if (_T_705) begin
                    if (_T_706) begin
                      if (_T_511) begin
                        if (_T_550) begin
                          Xstart_9 <= _GEN_105;
                        end else begin
                          Xstart_9 <= _T_546;
                        end
                      end else begin
                        Xstart_9 <= _T_546;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_10 <= 11'sh320;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_10 <= _T_372;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (_T_570) begin
                if (_T_511) begin
                  if (_T_577) begin
                    Xstart_10 <= _GEN_105;
                  end else begin
                    Xstart_10 <= _T_573;
                  end
                end else begin
                  Xstart_10 <= _T_573;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_11 <= 11'sh2a8;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_11 <= _T_375;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (_T_570) begin
                if (_T_511) begin
                  if (_T_595) begin
                    Xstart_11 <= _GEN_105;
                  end else begin
                    Xstart_11 <= _T_591;
                  end
                end else begin
                  Xstart_11 <= _T_591;
                end
              end else if (!(_T_627)) begin
                if (!(_T_684)) begin
                  if (_T_705) begin
                    if (_T_706) begin
                      if (_T_511) begin
                        if (_T_595) begin
                          Xstart_11 <= _GEN_105;
                        end else begin
                          Xstart_11 <= _T_591;
                        end
                      end else begin
                        Xstart_11 <= _T_591;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_12 <= 11'sh2ee;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_12 <= _T_378;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (_T_570) begin
                if (_T_511) begin
                  if (_T_613) begin
                    Xstart_12 <= _GEN_105;
                  end else begin
                    Xstart_12 <= _T_609;
                  end
                end else begin
                  Xstart_12 <= _T_609;
                end
              end else if (!(_T_627)) begin
                if (!(_T_684)) begin
                  if (_T_705) begin
                    if (_T_706) begin
                      if (_T_511) begin
                        if (_T_613) begin
                          Xstart_12 <= _GEN_105;
                        end else begin
                          Xstart_12 <= _T_609;
                        end
                      end else begin
                        Xstart_12 <= _T_609;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_13 <= 11'sh320;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_13 <= _T_381;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (_T_627) begin
                  if (_T_511) begin
                    if (_T_634) begin
                      Xstart_13 <= _GEN_105;
                    end else begin
                      Xstart_13 <= _T_630;
                    end
                  end else begin
                    Xstart_13 <= _T_630;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_14 <= 11'sh3d4;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_14 <= _T_384;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (_T_627) begin
                  if (_T_511) begin
                    if (_T_652) begin
                      Xstart_14 <= _GEN_105;
                    end else begin
                      Xstart_14 <= _T_648;
                    end
                  end else begin
                    Xstart_14 <= _T_648;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_15 <= 11'sh37a;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_15 <= _T_387;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (_T_627) begin
                  if (_T_511) begin
                    if (_T_670) begin
                      Xstart_15 <= _GEN_105;
                    end else begin
                      Xstart_15 <= _T_666;
                    end
                  end else begin
                    Xstart_15 <= _T_666;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_16 <= 11'sh258;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        Xstart_16 <= _T_390;
      end else if (!(_T_404)) begin
        if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (_T_684) begin
                    if (_T_688) begin
                      if (_T_691) begin
                        Xstart_16 <= _GEN_105;
                      end else begin
                        Xstart_16 <= _T_687;
                      end
                    end else begin
                      Xstart_16 <= _T_687;
                    end
                  end else if (_T_705) begin
                    if (_T_706) begin
                      if (_T_688) begin
                        if (_T_691) begin
                          Xstart_16 <= _GEN_105;
                        end else begin
                          Xstart_16 <= _T_687;
                        end
                      end else begin
                        Xstart_16 <= _T_687;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_17 <= 11'sh80;
    end else if (_T_341) begin
      Xstart_17 <= _T_288;
    end else if (_T_342) begin
      Xstart_17 <= _T_393;
    end else if (_T_404) begin
      Xstart_17 <= _T_288;
    end else if (_T_451) begin
      Xstart_17 <= _T_288;
    end else if (_T_486) begin
      Xstart_17 <= _T_288;
    end else if (_T_505) begin
      Xstart_17 <= _T_288;
    end else if (_T_570) begin
      Xstart_17 <= _T_288;
    end else if (_T_627) begin
      Xstart_17 <= _T_288;
    end else if (_T_684) begin
      Xstart_17 <= _T_288;
    end else if (_T_705) begin
      if (_T_830) begin
        if (_T_833) begin
          Xstart_17 <= _T_525;
        end else if (_T_825) begin
          Xstart_17 <= _T_828;
        end else begin
          Xstart_17 <= 11'sh1e0;
        end
      end else if (_T_825) begin
        Xstart_17 <= _T_828;
      end else begin
        Xstart_17 <= 11'sh1e0;
      end
    end else begin
      Xstart_17 <= _T_288;
    end
    if (reset) begin
      Xstart_18 <= 11'sh60;
    end else begin
      Xstart_18 <= _T_294;
    end
    if (reset) begin
      Xstart_19 <= 11'sh80;
    end else begin
      Xstart_19 <= _T_300;
    end
    if (reset) begin
      Xstart_20 <= 11'sh40;
    end else begin
      Xstart_20 <= _T_288;
    end
    if (reset) begin
      Xstart_21 <= 11'sh60;
    end else begin
      Xstart_21 <= _T_294;
    end
    if (reset) begin
      Xstart_22 <= 11'sh80;
    end else begin
      Xstart_22 <= _T_300;
    end
    if (reset) begin
      Xstart_23 <= 11'sh40;
    end else begin
      Xstart_23 <= _T_288;
    end
    if (reset) begin
      Xstart_24 <= 11'sh60;
    end else begin
      Xstart_24 <= _T_294;
    end
    if (reset) begin
      Xstart_25 <= 11'sh80;
    end else begin
      Xstart_25 <= _T_300;
    end
    if (reset) begin
      Xstart_26 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Xstart_26 <= 11'sh100;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_27 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Xstart_27 <= 11'sh120;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_28 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Xstart_28 <= 11'sh140;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_29 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Xstart_29 <= 11'sh160;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_30 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Xstart_30 <= 11'sh100;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_31 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Xstart_31 <= 11'sh120;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_32 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Xstart_32 <= 11'sh140;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_33 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Xstart_33 <= 11'sh160;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_41 <= 11'sh2bc;
    end else begin
      Xstart_41 <= Xstart_0;
    end
    if (reset) begin
      Xstart_42 <= 11'sh2bc;
    end else begin
      Xstart_42 <= Xstart_0;
    end
    if (reset) begin
      Xstart_43 <= 11'sh2bc;
    end else begin
      Xstart_43 <= Xstart_0;
    end
    if (reset) begin
      Xstart_44 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_44 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_45 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_45 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_46 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_46 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_47 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_47 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_48 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_48 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_49 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_49 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_50 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_50 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_51 <= 11'sh2bc;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              Xstart_51 <= 11'sh40;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_122 <= 11'sh2c0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1042) begin
                                  Xstart_122 <= _T_525;
                                end else begin
                                  Xstart_122 <= _T_1041;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_123 <= 11'sh2c0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1028) begin
                                  if (_T_1057) begin
                                    Xstart_123 <= _T_525;
                                  end else begin
                                    Xstart_123 <= _T_1056;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_124 <= 11'sh2c0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1029) begin
                                  if (_T_1070) begin
                                    Xstart_124 <= _T_525;
                                  end else begin
                                    Xstart_124 <= _T_1069;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_125 <= 11'sh2c0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_992) begin
                                Xstart_125 <= _T_525;
                              end else begin
                                Xstart_125 <= _T_991;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_126 <= 11'sh2c0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_978) begin
                                if (_T_1007) begin
                                  Xstart_126 <= _T_525;
                                end else begin
                                  Xstart_126 <= _T_1006;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Xstart_127 <= 11'sh2c0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_979) begin
                                if (_T_1020) begin
                                  Xstart_127 <= _T_525;
                                end else begin
                                  Xstart_127 <= _T_1019;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_0 <= 11'sh148;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (_T_862) begin
                          if (_T_863) begin
                            if (io_btnD) begin
                              if (_T_864) begin
                                Ystart_0 <= _T_867;
                              end
                            end else if (io_btnU) begin
                              if (_T_868) begin
                                Ystart_0 <= _T_871;
                              end
                            end
                          end
                        end else if (!(_T_886)) begin
                          if (_T_977) begin
                            if (die_10) begin
                              if (_T_1134) begin
                                Ystart_0 <= 11'she0;
                              end else if (die_9) begin
                                if (_T_1134) begin
                                  Ystart_0 <= 11'she0;
                                end else if (die_8) begin
                                  if (_T_1134) begin
                                    Ystart_0 <= 11'she0;
                                  end else if (die_7) begin
                                    if (_T_1134) begin
                                      Ystart_0 <= 11'she0;
                                    end else if (die_6) begin
                                      if (_T_1134) begin
                                        Ystart_0 <= 11'she0;
                                      end else if (die_5) begin
                                        if (_T_1134) begin
                                          Ystart_0 <= 11'she0;
                                        end else if (die_4) begin
                                          if (_T_1134) begin
                                            Ystart_0 <= 11'she0;
                                          end else if (die_3) begin
                                            if (_T_1134) begin
                                              Ystart_0 <= 11'she0;
                                            end else if (die_2) begin
                                              if (_T_1134) begin
                                                Ystart_0 <= 11'she0;
                                              end else if (die_1) begin
                                                if (_T_1134) begin
                                                  Ystart_0 <= 11'she0;
                                                end else if (die_0) begin
                                                  if (_T_1134) begin
                                                    Ystart_0 <= 11'she0;
                                                  end
                                                end
                                              end else if (die_0) begin
                                                if (_T_1134) begin
                                                  Ystart_0 <= 11'she0;
                                                end
                                              end
                                            end else if (die_1) begin
                                              if (_T_1134) begin
                                                Ystart_0 <= 11'she0;
                                              end else if (die_0) begin
                                                if (_T_1134) begin
                                                  Ystart_0 <= 11'she0;
                                                end
                                              end
                                            end else if (die_0) begin
                                              if (_T_1134) begin
                                                Ystart_0 <= 11'she0;
                                              end
                                            end
                                          end else if (die_2) begin
                                            if (_T_1134) begin
                                              Ystart_0 <= 11'she0;
                                            end else if (die_1) begin
                                              if (_T_1134) begin
                                                Ystart_0 <= 11'she0;
                                              end else begin
                                                Ystart_0 <= _GEN_1183;
                                              end
                                            end else begin
                                              Ystart_0 <= _GEN_1183;
                                            end
                                          end else if (die_1) begin
                                            if (_T_1134) begin
                                              Ystart_0 <= 11'she0;
                                            end else begin
                                              Ystart_0 <= _GEN_1183;
                                            end
                                          end else begin
                                            Ystart_0 <= _GEN_1183;
                                          end
                                        end else if (die_3) begin
                                          if (_T_1134) begin
                                            Ystart_0 <= 11'she0;
                                          end else if (die_2) begin
                                            if (_T_1134) begin
                                              Ystart_0 <= 11'she0;
                                            end else begin
                                              Ystart_0 <= _GEN_1193;
                                            end
                                          end else begin
                                            Ystart_0 <= _GEN_1193;
                                          end
                                        end else if (die_2) begin
                                          if (_T_1134) begin
                                            Ystart_0 <= 11'she0;
                                          end else begin
                                            Ystart_0 <= _GEN_1193;
                                          end
                                        end else begin
                                          Ystart_0 <= _GEN_1193;
                                        end
                                      end else if (die_4) begin
                                        if (_T_1134) begin
                                          Ystart_0 <= 11'she0;
                                        end else if (die_3) begin
                                          if (_T_1134) begin
                                            Ystart_0 <= 11'she0;
                                          end else begin
                                            Ystart_0 <= _GEN_1203;
                                          end
                                        end else begin
                                          Ystart_0 <= _GEN_1203;
                                        end
                                      end else if (die_3) begin
                                        if (_T_1134) begin
                                          Ystart_0 <= 11'she0;
                                        end else begin
                                          Ystart_0 <= _GEN_1203;
                                        end
                                      end else begin
                                        Ystart_0 <= _GEN_1203;
                                      end
                                    end else if (die_5) begin
                                      if (_T_1134) begin
                                        Ystart_0 <= 11'she0;
                                      end else if (die_4) begin
                                        if (_T_1134) begin
                                          Ystart_0 <= 11'she0;
                                        end else begin
                                          Ystart_0 <= _GEN_1213;
                                        end
                                      end else begin
                                        Ystart_0 <= _GEN_1213;
                                      end
                                    end else if (die_4) begin
                                      if (_T_1134) begin
                                        Ystart_0 <= 11'she0;
                                      end else begin
                                        Ystart_0 <= _GEN_1213;
                                      end
                                    end else begin
                                      Ystart_0 <= _GEN_1213;
                                    end
                                  end else if (die_6) begin
                                    if (_T_1134) begin
                                      Ystart_0 <= 11'she0;
                                    end else if (die_5) begin
                                      if (_T_1134) begin
                                        Ystart_0 <= 11'she0;
                                      end else begin
                                        Ystart_0 <= _GEN_1223;
                                      end
                                    end else begin
                                      Ystart_0 <= _GEN_1223;
                                    end
                                  end else if (die_5) begin
                                    if (_T_1134) begin
                                      Ystart_0 <= 11'she0;
                                    end else begin
                                      Ystart_0 <= _GEN_1223;
                                    end
                                  end else begin
                                    Ystart_0 <= _GEN_1223;
                                  end
                                end else if (die_7) begin
                                  if (_T_1134) begin
                                    Ystart_0 <= 11'she0;
                                  end else if (die_6) begin
                                    if (_T_1134) begin
                                      Ystart_0 <= 11'she0;
                                    end else begin
                                      Ystart_0 <= _GEN_1233;
                                    end
                                  end else begin
                                    Ystart_0 <= _GEN_1233;
                                  end
                                end else if (die_6) begin
                                  if (_T_1134) begin
                                    Ystart_0 <= 11'she0;
                                  end else begin
                                    Ystart_0 <= _GEN_1233;
                                  end
                                end else begin
                                  Ystart_0 <= _GEN_1233;
                                end
                              end else if (die_8) begin
                                if (_T_1134) begin
                                  Ystart_0 <= 11'she0;
                                end else if (die_7) begin
                                  if (_T_1134) begin
                                    Ystart_0 <= 11'she0;
                                  end else begin
                                    Ystart_0 <= _GEN_1243;
                                  end
                                end else begin
                                  Ystart_0 <= _GEN_1243;
                                end
                              end else if (die_7) begin
                                if (_T_1134) begin
                                  Ystart_0 <= 11'she0;
                                end else begin
                                  Ystart_0 <= _GEN_1243;
                                end
                              end else begin
                                Ystart_0 <= _GEN_1243;
                              end
                            end else if (die_9) begin
                              if (_T_1134) begin
                                Ystart_0 <= 11'she0;
                              end else if (die_8) begin
                                if (_T_1134) begin
                                  Ystart_0 <= 11'she0;
                                end else begin
                                  Ystart_0 <= _GEN_1253;
                                end
                              end else begin
                                Ystart_0 <= _GEN_1253;
                              end
                            end else if (die_8) begin
                              if (_T_1134) begin
                                Ystart_0 <= 11'she0;
                              end else begin
                                Ystart_0 <= _GEN_1253;
                              end
                            end else begin
                              Ystart_0 <= _GEN_1253;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_1 <= 11'sh148;
    end else begin
      Ystart_1 <= Ystart_0;
    end
    if (reset) begin
      Ystart_2 <= 11'sh64;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (!(_T_909)) begin
                                if (!(_T_924)) begin
                                  if (shotPop_0) begin
                                    if (shotLoad) begin
                                      Ystart_2 <= _T_945;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_3 <= 11'sh96;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (!(_T_909)) begin
                                if (!(_T_924)) begin
                                  if (!(shotPop_0)) begin
                                    if (shotPop_1) begin
                                      if (shotLoad) begin
                                        Ystart_3 <= _T_958;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_4 <= 11'sh64;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (!(_T_909)) begin
                                if (!(_T_924)) begin
                                  if (!(shotPop_0)) begin
                                    if (!(shotPop_1)) begin
                                      if (shotPop_2) begin
                                        if (shotLoad) begin
                                          Ystart_4 <= _T_971;
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_5 <= 11'sh64;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (_T_909) begin
                                if (shotPop_3) begin
                                  if (shotLoad) begin
                                    Ystart_5 <= _T_917;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_6 <= 11'sh64;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (!(_T_909)) begin
                                if (_T_924) begin
                                  if (shotPop_4) begin
                                    if (shotLoad) begin
                                      Ystart_6 <= _T_932;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_7 <= 11'sh64;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (_T_505) begin
                if (_T_507) begin
                  if (_T_511) begin
                    if (_T_514) begin
                      if (_T_501) begin
                        Ystart_7 <= _T_521;
                      end else begin
                        Ystart_7 <= {{1{Randomizer_io_out[9]}},Randomizer_io_out};
                      end
                    end
                  end
                end
              end else if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (_T_705) begin
                      if (_T_706) begin
                        if (_T_511) begin
                          if (_T_514) begin
                            if (_T_501) begin
                              Ystart_7 <= _T_720;
                            end else begin
                              Ystart_7 <= {{1{Randomizer_20_io_out[9]}},Randomizer_20_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_8 <= 11'sh7d;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (_T_505) begin
                if (_T_507) begin
                  if (_T_511) begin
                    if (_T_532) begin
                      if (_T_501) begin
                        Ystart_8 <= _T_539;
                      end else begin
                        Ystart_8 <= {{1{Randomizer_2_io_out[9]}},Randomizer_2_io_out};
                      end
                    end
                  end
                end
              end else if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (_T_705) begin
                      if (_T_706) begin
                        if (_T_511) begin
                          if (_T_532) begin
                            if (_T_501) begin
                              Ystart_8 <= _T_738;
                            end else begin
                              Ystart_8 <= {{1{Randomizer_22_io_out[9]}},Randomizer_22_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_9 <= 11'sh96;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (_T_505) begin
                if (_T_507) begin
                  if (_T_511) begin
                    if (_T_550) begin
                      if (_T_501) begin
                        Ystart_9 <= _T_557;
                      end else begin
                        Ystart_9 <= {{1{Randomizer_4_io_out[9]}},Randomizer_4_io_out};
                      end
                    end
                  end
                end
              end else if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (_T_705) begin
                      if (_T_706) begin
                        if (_T_511) begin
                          if (_T_550) begin
                            if (_T_501) begin
                              Ystart_9 <= _T_756;
                            end else begin
                              Ystart_9 <= {{1{Randomizer_24_io_out[9]}},Randomizer_24_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_10 <= 11'shaa;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (_T_570) begin
                  if (_T_511) begin
                    if (_T_577) begin
                      if (_T_501) begin
                        Ystart_10 <= _T_584;
                      end else begin
                        Ystart_10 <= {{1{Randomizer_6_io_out[9]}},Randomizer_6_io_out};
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_11 <= 11'shb4;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (_T_570) begin
                  if (_T_511) begin
                    if (_T_595) begin
                      if (_T_501) begin
                        Ystart_11 <= _T_602;
                      end else begin
                        Ystart_11 <= {{1{Randomizer_8_io_out[9]}},Randomizer_8_io_out};
                      end
                    end
                  end
                end else if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (_T_705) begin
                      if (_T_706) begin
                        if (_T_511) begin
                          if (_T_595) begin
                            if (_T_501) begin
                              Ystart_11 <= _T_774;
                            end else begin
                              Ystart_11 <= {{1{Randomizer_26_io_out[9]}},Randomizer_26_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_12 <= 11'shc8;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (_T_570) begin
                  if (_T_511) begin
                    if (_T_613) begin
                      if (_T_501) begin
                        Ystart_12 <= _T_620;
                      end else begin
                        Ystart_12 <= {{1{Randomizer_10_io_out[9]}},Randomizer_10_io_out};
                      end
                    end
                  end
                end else if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (_T_705) begin
                      if (_T_706) begin
                        if (_T_511) begin
                          if (_T_613) begin
                            if (_T_501) begin
                              Ystart_12 <= _T_792;
                            end else begin
                              Ystart_12 <= {{1{Randomizer_28_io_out[9]}},Randomizer_28_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_13 <= 11'shfa;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (_T_627) begin
                    if (_T_511) begin
                      if (_T_634) begin
                        if (_T_501) begin
                          Ystart_13 <= _T_641;
                        end else begin
                          Ystart_13 <= {{1{Randomizer_12_io_out[9]}},Randomizer_12_io_out};
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_14 <= 11'sh12c;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (_T_627) begin
                    if (_T_511) begin
                      if (_T_652) begin
                        if (_T_501) begin
                          Ystart_14 <= _T_659;
                        end else begin
                          Ystart_14 <= {{1{Randomizer_14_io_out[9]}},Randomizer_14_io_out};
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_15 <= 11'sh14c;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (_T_627) begin
                    if (_T_511) begin
                      if (_T_670) begin
                        if (_T_501) begin
                          Ystart_15 <= _T_677;
                        end else begin
                          Ystart_15 <= {{1{Randomizer_16_io_out[9]}},Randomizer_16_io_out};
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_16 <= 11'shc8;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (_T_684) begin
                      if (_T_688) begin
                        if (_T_691) begin
                          if (_T_501) begin
                            Ystart_16 <= _T_698;
                          end else begin
                            Ystart_16 <= {{1{Randomizer_18_io_out[9]}},Randomizer_18_io_out};
                          end
                        end
                      end
                    end else if (_T_705) begin
                      if (_T_706) begin
                        if (_T_688) begin
                          if (_T_691) begin
                            if (_T_501) begin
                              Ystart_16 <= _T_810;
                            end else begin
                              Ystart_16 <= {{1{Randomizer_30_io_out[9]}},Randomizer_30_io_out};
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_17 <= 11'sh80;
    end else if (_T_341) begin
      Ystart_17 <= _T_291;
    end else if (_T_342) begin
      Ystart_17 <= _T_291;
    end else if (_T_404) begin
      Ystart_17 <= _T_291;
    end else if (_T_451) begin
      Ystart_17 <= _T_291;
    end else if (_T_486) begin
      Ystart_17 <= _T_291;
    end else if (_T_505) begin
      Ystart_17 <= _T_291;
    end else if (_T_570) begin
      Ystart_17 <= _T_291;
    end else if (_T_627) begin
      Ystart_17 <= _T_291;
    end else if (_T_684) begin
      Ystart_17 <= _T_291;
    end else if (_T_705) begin
      if (_T_830) begin
        if (_T_833) begin
          Ystart_17 <= {{1{_T_845[9]}},_T_845};
        end else begin
          Ystart_17 <= _T_824;
        end
      end else begin
        Ystart_17 <= _T_824;
      end
    end else begin
      Ystart_17 <= _T_291;
    end
    if (reset) begin
      Ystart_18 <= 11'sh40;
    end else begin
      Ystart_18 <= _T_291;
    end
    if (reset) begin
      Ystart_19 <= 11'sh40;
    end else begin
      Ystart_19 <= _T_291;
    end
    if (reset) begin
      Ystart_20 <= 11'sh60;
    end else begin
      Ystart_20 <= _T_309;
    end
    if (reset) begin
      Ystart_21 <= 11'sh60;
    end else begin
      Ystart_21 <= _T_309;
    end
    if (reset) begin
      Ystart_22 <= 11'sh60;
    end else begin
      Ystart_22 <= _T_309;
    end
    if (reset) begin
      Ystart_23 <= 11'sh80;
    end else begin
      Ystart_23 <= _T_327;
    end
    if (reset) begin
      Ystart_24 <= 11'sh80;
    end else begin
      Ystart_24 <= _T_327;
    end
    if (reset) begin
      Ystart_25 <= 11'sh80;
    end else begin
      Ystart_25 <= _T_327;
    end
    if (reset) begin
      Ystart_26 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Ystart_26 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_27 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Ystart_27 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_28 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Ystart_28 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_29 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_281) begin
                                Ystart_29 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_30 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Ystart_30 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_31 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Ystart_31 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_32 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Ystart_32 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_33 <= 11'sh20;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_500) begin
                                Ystart_33 <= 11'she0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_41 <= 11'sh20;
    end else begin
      Ystart_41 <= Ystart_0;
    end
    if (reset) begin
      Ystart_42 <= 11'sh20;
    end else begin
      Ystart_42 <= Ystart_0;
    end
    if (reset) begin
      Ystart_43 <= 11'sh20;
    end else begin
      Ystart_43 <= Ystart_0;
    end
    if (reset) begin
      Ystart_122 <= 11'sh96;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1042) begin
                                  Ystart_122 <= {{1{Randomizer_41_io_out[9]}},Randomizer_41_io_out};
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_123 <= 11'shfa;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1028) begin
                                  if (_T_1057) begin
                                    Ystart_123 <= {{1{Randomizer_43_io_out[9]}},Randomizer_43_io_out};
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_124 <= 11'sh140;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1029) begin
                                  if (_T_1070) begin
                                    Ystart_124 <= {{1{Randomizer_45_io_out[9]}},Randomizer_45_io_out};
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_125 <= 11'shd2;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_992) begin
                                Ystart_125 <= {{1{Randomizer_34_io_out[9]}},Randomizer_34_io_out};
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_126 <= 11'sh64;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_978) begin
                                if (_T_1007) begin
                                  Ystart_126 <= {{1{Randomizer_36_io_out[9]}},Randomizer_36_io_out};
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      Ystart_127 <= 11'sh12c;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_979) begin
                                if (_T_1020) begin
                                  Ystart_127 <= {{1{Randomizer_38_io_out[9]}},Randomizer_38_io_out};
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    spriteVisibleReg_0 <= reset | _GEN_0;
    spriteVisibleReg_1 <= reset | _GEN_1;
    spriteVisibleReg_2 <= reset | _GEN_4158;
    spriteVisibleReg_3 <= reset | _GEN_4161;
    spriteVisibleReg_4 <= reset | _GEN_4164;
    spriteVisibleReg_5 <= reset | _GEN_4167;
    spriteVisibleReg_6 <= reset | _GEN_4170;
    if (reset) begin
      spriteVisibleReg_7 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_7 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_505) begin
      if (_T_507) begin
        if (kill_0_4) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_3) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_2) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_1) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_0) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_7 <= _GEN_108;
        end else begin
          spriteVisibleReg_7 <= _GEN_9;
        end
      end else begin
        spriteVisibleReg_7 <= _GEN_9;
      end
    end else if (_T_570) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_627) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_684) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_0_4) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_3) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_2) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_1) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (kill_0_0) begin
          spriteVisibleReg_7 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_7 <= _GEN_108;
        end else begin
          spriteVisibleReg_7 <= _GEN_9;
        end
      end else begin
        spriteVisibleReg_7 <= _GEN_9;
      end
    end else if (_T_862) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_886) begin
      spriteVisibleReg_7 <= _GEN_9;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_7 <= 1'h0;
      end else begin
        spriteVisibleReg_7 <= _GEN_9;
      end
    end else begin
      spriteVisibleReg_7 <= _GEN_9;
    end
    if (reset) begin
      spriteVisibleReg_8 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_8 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_505) begin
      if (_T_507) begin
        if (kill_1_4) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_3) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_2) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_1) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_0) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_8 <= _GEN_158;
        end else begin
          spriteVisibleReg_8 <= _GEN_11;
        end
      end else begin
        spriteVisibleReg_8 <= _GEN_11;
      end
    end else if (_T_570) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_627) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_684) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_1_4) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_3) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_2) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_1) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (kill_1_0) begin
          spriteVisibleReg_8 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_8 <= _GEN_158;
        end else begin
          spriteVisibleReg_8 <= _GEN_11;
        end
      end else begin
        spriteVisibleReg_8 <= _GEN_11;
      end
    end else if (_T_862) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_886) begin
      spriteVisibleReg_8 <= _GEN_11;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_8 <= 1'h0;
      end else begin
        spriteVisibleReg_8 <= _GEN_11;
      end
    end else begin
      spriteVisibleReg_8 <= _GEN_11;
    end
    if (reset) begin
      spriteVisibleReg_9 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_9 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_505) begin
      if (_T_507) begin
        if (kill_2_4) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_3) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_2) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_1) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_0) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_9 <= _GEN_208;
        end else begin
          spriteVisibleReg_9 <= _GEN_13;
        end
      end else begin
        spriteVisibleReg_9 <= _GEN_13;
      end
    end else if (_T_570) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_627) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_684) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_2_4) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_3) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_2) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_1) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (kill_2_0) begin
          spriteVisibleReg_9 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_9 <= _GEN_208;
        end else begin
          spriteVisibleReg_9 <= _GEN_13;
        end
      end else begin
        spriteVisibleReg_9 <= _GEN_13;
      end
    end else if (_T_862) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_886) begin
      spriteVisibleReg_9 <= _GEN_13;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_9 <= 1'h0;
      end else begin
        spriteVisibleReg_9 <= _GEN_13;
      end
    end else begin
      spriteVisibleReg_9 <= _GEN_13;
    end
    if (reset) begin
      spriteVisibleReg_10 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_10 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_505) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_570) begin
      if (kill_3_4) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_3) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_2) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_1) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (kill_3_0) begin
        spriteVisibleReg_10 <= 1'h0;
      end else if (_T_511) begin
        spriteVisibleReg_10 <= _GEN_286;
      end else begin
        spriteVisibleReg_10 <= _GEN_15;
      end
    end else if (_T_627) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_684) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_705) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_862) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_886) begin
      spriteVisibleReg_10 <= _GEN_15;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_10 <= 1'h0;
      end else begin
        spriteVisibleReg_10 <= _GEN_15;
      end
    end else begin
      spriteVisibleReg_10 <= _GEN_15;
    end
    if (reset) begin
      spriteVisibleReg_11 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_11 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_505) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_570) begin
      if (kill_4_4) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_3) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_2) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_1) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (kill_4_0) begin
        spriteVisibleReg_11 <= 1'h0;
      end else if (_T_511) begin
        spriteVisibleReg_11 <= _GEN_336;
      end else begin
        spriteVisibleReg_11 <= _GEN_17;
      end
    end else if (_T_627) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_684) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_4_4) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_3) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_2) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_1) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (kill_4_0) begin
          spriteVisibleReg_11 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_11 <= _GEN_336;
        end else begin
          spriteVisibleReg_11 <= _GEN_17;
        end
      end else begin
        spriteVisibleReg_11 <= _GEN_17;
      end
    end else if (_T_862) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_886) begin
      spriteVisibleReg_11 <= _GEN_17;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_11 <= 1'h0;
      end else begin
        spriteVisibleReg_11 <= _GEN_17;
      end
    end else begin
      spriteVisibleReg_11 <= _GEN_17;
    end
    if (reset) begin
      spriteVisibleReg_12 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_12 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_505) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_570) begin
      if (kill_5_4) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_3) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_2) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_1) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (kill_5_0) begin
        spriteVisibleReg_12 <= 1'h0;
      end else if (_T_511) begin
        spriteVisibleReg_12 <= _GEN_386;
      end else begin
        spriteVisibleReg_12 <= _GEN_19;
      end
    end else if (_T_627) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_684) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_5_4) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_3) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_2) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_1) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (kill_5_0) begin
          spriteVisibleReg_12 <= 1'h0;
        end else if (_T_511) begin
          spriteVisibleReg_12 <= _GEN_386;
        end else begin
          spriteVisibleReg_12 <= _GEN_19;
        end
      end else begin
        spriteVisibleReg_12 <= _GEN_19;
      end
    end else if (_T_862) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_886) begin
      spriteVisibleReg_12 <= _GEN_19;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_12 <= 1'h0;
      end else begin
        spriteVisibleReg_12 <= _GEN_19;
      end
    end else begin
      spriteVisibleReg_12 <= _GEN_19;
    end
    if (reset) begin
      spriteVisibleReg_13 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_13 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_505) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_570) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_627) begin
      if (kill_6_4) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_3) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_2) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_1) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (kill_6_0) begin
        spriteVisibleReg_13 <= 1'h0;
      end else if (_T_511) begin
        spriteVisibleReg_13 <= _GEN_436;
      end else begin
        spriteVisibleReg_13 <= _GEN_21;
      end
    end else if (_T_684) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_705) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_862) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_886) begin
      spriteVisibleReg_13 <= _GEN_21;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_13 <= 1'h0;
      end else begin
        spriteVisibleReg_13 <= _GEN_21;
      end
    end else begin
      spriteVisibleReg_13 <= _GEN_21;
    end
    if (reset) begin
      spriteVisibleReg_14 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_14 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_505) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_570) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_627) begin
      if (kill_7_4) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_3) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_2) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_1) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (kill_7_0) begin
        spriteVisibleReg_14 <= 1'h0;
      end else if (_T_511) begin
        spriteVisibleReg_14 <= _GEN_486;
      end else begin
        spriteVisibleReg_14 <= _GEN_23;
      end
    end else if (_T_684) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_705) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_862) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_886) begin
      spriteVisibleReg_14 <= _GEN_23;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_14 <= 1'h0;
      end else begin
        spriteVisibleReg_14 <= _GEN_23;
      end
    end else begin
      spriteVisibleReg_14 <= _GEN_23;
    end
    if (reset) begin
      spriteVisibleReg_15 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_15 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_505) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_570) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_627) begin
      if (kill_8_4) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_3) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_2) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_1) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (kill_8_0) begin
        spriteVisibleReg_15 <= 1'h0;
      end else if (_T_511) begin
        spriteVisibleReg_15 <= _GEN_536;
      end else begin
        spriteVisibleReg_15 <= _GEN_25;
      end
    end else if (_T_684) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_705) begin
      spriteVisibleReg_15 <= 1'h0;
    end else if (_T_862) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_886) begin
      spriteVisibleReg_15 <= _GEN_25;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_15 <= 1'h0;
      end else begin
        spriteVisibleReg_15 <= _GEN_25;
      end
    end else begin
      spriteVisibleReg_15 <= _GEN_25;
    end
    if (reset) begin
      spriteVisibleReg_16 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_16 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_505) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_570) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_627) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_684) begin
      if (kill_9_3) begin
        spriteVisibleReg_16 <= 1'h0;
      end else if (_T_688) begin
        spriteVisibleReg_16 <= _GEN_586;
      end else begin
        spriteVisibleReg_16 <= _GEN_27;
      end
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_9_3) begin
          spriteVisibleReg_16 <= 1'h0;
        end else if (_T_688) begin
          spriteVisibleReg_16 <= _GEN_586;
        end else begin
          spriteVisibleReg_16 <= _GEN_27;
        end
      end else begin
        spriteVisibleReg_16 <= _GEN_27;
      end
    end else if (_T_862) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_886) begin
      spriteVisibleReg_16 <= _GEN_27;
    end else if (_T_977) begin
      if (_T_1085) begin
        spriteVisibleReg_16 <= 1'h0;
      end else begin
        spriteVisibleReg_16 <= _GEN_27;
      end
    end else begin
      spriteVisibleReg_16 <= _GEN_27;
    end
    if (reset) begin
      spriteVisibleReg_17 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        spriteVisibleReg_17 <= 1'h0;
      end
    end else if (_T_486) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_505) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_570) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_627) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_684) begin
      spriteVisibleReg_17 <= _GEN_29;
    end else if (_T_705) begin
      if (_T_500) begin
        spriteVisibleReg_17 <= 1'h0;
      end else if (_T_830) begin
        spriteVisibleReg_17 <= _GEN_827;
      end else begin
        spriteVisibleReg_17 <= _GEN_29;
      end
    end else begin
      spriteVisibleReg_17 <= _GEN_29;
    end
    spriteVisibleReg_18 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_19 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_20 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_21 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_22 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_23 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_24 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_25 <= reset | spriteVisibleReg_17;
    spriteVisibleReg_26 <= reset | _GEN_4318;
    spriteVisibleReg_27 <= reset | _GEN_4324;
    spriteVisibleReg_28 <= reset | _GEN_4330;
    spriteVisibleReg_29 <= reset | _GEN_4336;
    spriteVisibleReg_30 <= reset | _GEN_4321;
    spriteVisibleReg_31 <= reset | _GEN_4327;
    spriteVisibleReg_32 <= reset | _GEN_4333;
    spriteVisibleReg_33 <= reset | _GEN_4339;
    spriteVisibleReg_41 <= reset | _GEN_4;
    spriteVisibleReg_42 <= reset | _GEN_5;
    spriteVisibleReg_43 <= reset | _GEN_6;
    spriteVisibleReg_44 <= reset | _GEN_4354;
    spriteVisibleReg_45 <= reset | _GEN_4357;
    spriteVisibleReg_46 <= reset | _GEN_4360;
    spriteVisibleReg_47 <= reset | _GEN_4363;
    spriteVisibleReg_48 <= reset | _GEN_4366;
    spriteVisibleReg_49 <= reset | _GEN_4369;
    spriteVisibleReg_50 <= reset | _GEN_4372;
    spriteVisibleReg_51 <= reset | _GEN_4375;
    spriteVisibleReg_55 <= reset | _GEN_4352;
    spriteVisibleReg_56 <= reset | _GEN_4348;
    spriteVisibleReg_57 <= reset | _GEN_4344;
    spriteVisibleReg_61 <= reset | _GEN_4345;
    spriteVisibleReg_62 <= reset | _GEN_4349;
    spriteVisibleReg_63 <= reset | _GEN_4353;
    spriteVisibleReg_64 <= reset | _GEN_4351;
    spriteVisibleReg_65 <= reset | _GEN_4347;
    spriteVisibleReg_66 <= reset | _GEN_4343;
    spriteVisibleReg_70 <= reset | _GEN_4350;
    spriteVisibleReg_71 <= reset | _GEN_4346;
    spriteVisibleReg_72 <= reset | _GEN_4342;
    if (reset) begin
      spriteFlipVerticalReg_122 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1042) begin
                                  spriteFlipVerticalReg_122 <= _T_1047;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_123 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1028) begin
                                  if (_T_1057) begin
                                    spriteFlipVerticalReg_123 <= _T_1062;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_124 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1027) begin
                                if (_T_1029) begin
                                  if (_T_1070) begin
                                    spriteFlipVerticalReg_124 <= _T_1075;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_125 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_992) begin
                                spriteFlipVerticalReg_125 <= _T_997;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_126 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_978) begin
                                if (_T_1007) begin
                                  spriteFlipVerticalReg_126 <= _T_1012;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spriteFlipVerticalReg_127 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_979) begin
                                if (_T_1020) begin
                                  spriteFlipVerticalReg_127 <= _T_1025;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btnCReg <= io_btnC;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              btnCReg <= io_btnC;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      viewX <= 10'h0;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        if (_T_395) begin
          viewX <= _T_401;
        end else begin
          viewX <= _T_345;
        end
      end
    end
    if (reset) begin
      stateReg <= 4'h0;
    end else if (_T_341) begin
      if (io_newFrame) begin
        stateReg <= 4'h1;
      end
    end else if (_T_342) begin
      if (levelCng) begin
        stateReg <= 4'h2;
      end else begin
        stateReg <= 4'h5;
      end
    end else if (_T_404) begin
      if (_T_437) begin
        if (_T_408) begin
          stateReg <= 4'h2;
        end else if (_T_423) begin
          if (_T_408) begin
            stateReg <= 4'h2;
          end else if (_T_406) begin
            if (_T_407) begin
              if (_T_408) begin
                stateReg <= 4'h2;
              end else begin
                stateReg <= 4'h3;
              end
            end else begin
              stateReg <= 4'h3;
            end
          end else begin
            stateReg <= 4'h3;
          end
        end else if (_T_406) begin
          if (_T_407) begin
            if (_T_408) begin
              stateReg <= 4'h2;
            end else begin
              stateReg <= 4'h3;
            end
          end else begin
            stateReg <= 4'h3;
          end
        end else begin
          stateReg <= 4'h3;
        end
      end else if (_T_423) begin
        if (_T_408) begin
          stateReg <= 4'h2;
        end else if (_T_406) begin
          if (_T_407) begin
            if (_T_408) begin
              stateReg <= 4'h2;
            end else begin
              stateReg <= 4'h3;
            end
          end else begin
            stateReg <= 4'h3;
          end
        end else begin
          stateReg <= 4'h3;
        end
      end else if (_T_406) begin
        if (_T_407) begin
          if (_T_408) begin
            stateReg <= 4'h2;
          end else begin
            stateReg <= 4'h3;
          end
        end else begin
          stateReg <= 4'h3;
        end
      end else begin
        stateReg <= 4'h3;
      end
    end else if (_T_451) begin
      if (_T_437) begin
        if (_T_408) begin
          stateReg <= 4'h3;
        end else if (_T_423) begin
          if (_T_408) begin
            stateReg <= 4'h3;
          end else begin
            stateReg <= 4'h4;
          end
        end else begin
          stateReg <= 4'h4;
        end
      end else if (_T_423) begin
        if (_T_408) begin
          stateReg <= 4'h3;
        end else begin
          stateReg <= 4'h4;
        end
      end else begin
        stateReg <= 4'h4;
      end
    end else if (_T_486) begin
      if (_T_408) begin
        stateReg <= 4'h4;
      end else if (_T_500) begin
        stateReg <= 4'ha;
      end else if (_T_503) begin
        stateReg <= 4'h9;
      end else begin
        stateReg <= 4'h5;
      end
    end else if (_T_505) begin
      if (_T_507) begin
        if (_T_562) begin
          if (_T_565) begin
            stateReg <= 4'h9;
          end else begin
            stateReg <= 4'h6;
          end
        end else begin
          stateReg <= 4'ha;
        end
      end else if (_T_502) begin
        stateReg <= 4'h9;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_570) begin
      if (_T_625) begin
        stateReg <= 4'h7;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_627) begin
      if (_T_682) begin
        stateReg <= 4'h8;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_684) begin
      if (_T_501) begin
        stateReg <= 4'h9;
      end else begin
        stateReg <= 4'ha;
      end
    end else if (_T_705) begin
      stateReg <= 4'ha;
    end else if (_T_862) begin
      if (_T_863) begin
        stateReg <= 4'hb;
      end else begin
        stateReg <= 4'hc;
      end
    end else if (_T_886) begin
      stateReg <= 4'hc;
    end else if (_T_977) begin
      stateReg <= 4'hd;
    end else if (_T_1455) begin
      stateReg <= 4'h0;
    end
    if (reset) begin
      shotCnt <= 10'shf;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (!(_T_909)) begin
                                if (!(_T_924)) begin
                                  if (shotPop_0) begin
                                    if (_T_919) begin
                                      shotCnt <= _T_950;
                                    end
                                  end else if (shotPop_1) begin
                                    if (_T_919) begin
                                      shotCnt <= _T_950;
                                    end
                                  end else if (shotPop_2) begin
                                    if (_T_919) begin
                                      shotCnt <= _T_950;
                                    end
                                  end
                                end
                              end
                            end
                          end else if (_T_977) begin
                            if (io_sw_0) begin
                              shotCnt <= 10'shf;
                            end else if (_T_1088) begin
                              if (_T_1099) begin
                                shotCnt <= 10'shf;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      shotLoad <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (_T_909) begin
                                if (shotPop_3) begin
                                  if (_T_919) begin
                                    shotLoad <= 1'h0;
                                  end else begin
                                    shotLoad <= _GEN_887;
                                  end
                                end
                              end else if (_T_924) begin
                                if (shotPop_4) begin
                                  if (_T_919) begin
                                    shotLoad <= 1'h0;
                                  end else begin
                                    shotLoad <= _GEN_902;
                                  end
                                end
                              end else if (shotPop_0) begin
                                if (_T_919) begin
                                  shotLoad <= 1'h0;
                                end else begin
                                  shotLoad <= _GEN_917;
                                end
                              end else if (shotPop_1) begin
                                if (_T_919) begin
                                  shotLoad <= 1'h0;
                                end else begin
                                  shotLoad <= _GEN_917;
                                end
                              end else if (shotPop_2) begin
                                if (_T_919) begin
                                  shotLoad <= 1'h0;
                                end else begin
                                  shotLoad <= _GEN_917;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      shotCntBig <= 3'sh3;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (_T_909) begin
                                if (shotPop_3) begin
                                  if (_T_919) begin
                                    shotCntBig <= _T_922;
                                  end
                                end
                              end
                            end
                          end else if (_T_977) begin
                            if (io_sw_0) begin
                              shotCntBig <= 3'sh3;
                            end else if (_T_1088) begin
                              if (_T_1099) begin
                                shotCntBig <= 3'sh3;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      shotCntFast <= 3'sh3;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (_T_886) begin
                            if (_T_863) begin
                              if (!(_T_909)) begin
                                if (_T_924) begin
                                  if (shotPop_4) begin
                                    if (_T_919) begin
                                      shotCntFast <= _T_937;
                                    end
                                  end
                                end
                              end
                            end
                          end else if (_T_977) begin
                            if (io_sw_0) begin
                              shotCntFast <= 3'sh3;
                            end else if (_T_1088) begin
                              if (_T_1099) begin
                                shotCntFast <= 3'sh3;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    shotPop_0 <= reset | _GEN_4157;
    shotPop_1 <= reset | _GEN_4160;
    shotPop_2 <= reset | _GEN_4163;
    shotPop_3 <= reset | _GEN_4166;
    shotPop_4 <= reset | _GEN_4169;
    shotInteract_0 <= reset | _GEN_4156;
    shotInteract_1 <= reset | _GEN_4159;
    shotInteract_2 <= reset | _GEN_4162;
    shotInteract_3 <= reset | _GEN_4165;
    shotInteract_4 <= reset | _GEN_4168;
    if (reset) begin
      astInteract_0 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_0 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_505) begin
      if (_T_507) begin
        if (kill_0_4) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_3) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_2) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_1) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_0) begin
          astInteract_0 <= 1'h0;
        end else if (_T_511) begin
          astInteract_0 <= _GEN_107;
        end else begin
          astInteract_0 <= _GEN_8;
        end
      end else begin
        astInteract_0 <= _GEN_8;
      end
    end else if (_T_570) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_627) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_684) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_0_4) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_3) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_2) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_1) begin
          astInteract_0 <= 1'h0;
        end else if (kill_0_0) begin
          astInteract_0 <= 1'h0;
        end else if (_T_511) begin
          astInteract_0 <= _GEN_107;
        end else begin
          astInteract_0 <= _GEN_8;
        end
      end else begin
        astInteract_0 <= _GEN_8;
      end
    end else if (_T_862) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_886) begin
      astInteract_0 <= _GEN_8;
    end else if (_T_977) begin
      if (die_0) begin
        if (_T_1136) begin
          astInteract_0 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_0 <= 1'h0;
        end else begin
          astInteract_0 <= _GEN_8;
        end
      end else if (_T_1085) begin
        astInteract_0 <= 1'h0;
      end else begin
        astInteract_0 <= _GEN_8;
      end
    end else begin
      astInteract_0 <= _GEN_8;
    end
    if (reset) begin
      astInteract_1 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_1 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_505) begin
      if (_T_507) begin
        if (kill_1_4) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_3) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_2) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_1) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_0) begin
          astInteract_1 <= 1'h0;
        end else if (_T_511) begin
          astInteract_1 <= _GEN_157;
        end else begin
          astInteract_1 <= _GEN_10;
        end
      end else begin
        astInteract_1 <= _GEN_10;
      end
    end else if (_T_570) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_627) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_684) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_1_4) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_3) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_2) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_1) begin
          astInteract_1 <= 1'h0;
        end else if (kill_1_0) begin
          astInteract_1 <= 1'h0;
        end else if (_T_511) begin
          astInteract_1 <= _GEN_157;
        end else begin
          astInteract_1 <= _GEN_10;
        end
      end else begin
        astInteract_1 <= _GEN_10;
      end
    end else if (_T_862) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_886) begin
      astInteract_1 <= _GEN_10;
    end else if (_T_977) begin
      if (die_1) begin
        if (_T_1136) begin
          astInteract_1 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_1 <= 1'h0;
        end else begin
          astInteract_1 <= _GEN_10;
        end
      end else if (_T_1085) begin
        astInteract_1 <= 1'h0;
      end else begin
        astInteract_1 <= _GEN_10;
      end
    end else begin
      astInteract_1 <= _GEN_10;
    end
    if (reset) begin
      astInteract_2 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_2 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_505) begin
      if (_T_507) begin
        if (kill_2_4) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_3) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_2) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_1) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_0) begin
          astInteract_2 <= 1'h0;
        end else if (_T_511) begin
          astInteract_2 <= _GEN_207;
        end else begin
          astInteract_2 <= _GEN_12;
        end
      end else begin
        astInteract_2 <= _GEN_12;
      end
    end else if (_T_570) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_627) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_684) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_2_4) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_3) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_2) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_1) begin
          astInteract_2 <= 1'h0;
        end else if (kill_2_0) begin
          astInteract_2 <= 1'h0;
        end else if (_T_511) begin
          astInteract_2 <= _GEN_207;
        end else begin
          astInteract_2 <= _GEN_12;
        end
      end else begin
        astInteract_2 <= _GEN_12;
      end
    end else if (_T_862) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_886) begin
      astInteract_2 <= _GEN_12;
    end else if (_T_977) begin
      if (die_2) begin
        if (_T_1136) begin
          astInteract_2 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_2 <= 1'h0;
        end else begin
          astInteract_2 <= _GEN_12;
        end
      end else if (_T_1085) begin
        astInteract_2 <= 1'h0;
      end else begin
        astInteract_2 <= _GEN_12;
      end
    end else begin
      astInteract_2 <= _GEN_12;
    end
    if (reset) begin
      astInteract_3 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_3 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_505) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_570) begin
      if (kill_3_4) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_3) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_2) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_1) begin
        astInteract_3 <= 1'h0;
      end else if (kill_3_0) begin
        astInteract_3 <= 1'h0;
      end else if (_T_511) begin
        astInteract_3 <= _GEN_285;
      end else begin
        astInteract_3 <= _GEN_14;
      end
    end else if (_T_627) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_684) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_705) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_862) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_886) begin
      astInteract_3 <= _GEN_14;
    end else if (_T_977) begin
      if (die_3) begin
        if (_T_1136) begin
          astInteract_3 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_3 <= 1'h0;
        end else begin
          astInteract_3 <= _GEN_14;
        end
      end else if (_T_1085) begin
        astInteract_3 <= 1'h0;
      end else begin
        astInteract_3 <= _GEN_14;
      end
    end else begin
      astInteract_3 <= _GEN_14;
    end
    if (reset) begin
      astInteract_4 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_4 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_505) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_570) begin
      if (kill_4_4) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_3) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_2) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_1) begin
        astInteract_4 <= 1'h0;
      end else if (kill_4_0) begin
        astInteract_4 <= 1'h0;
      end else if (_T_511) begin
        astInteract_4 <= _GEN_335;
      end else begin
        astInteract_4 <= _GEN_16;
      end
    end else if (_T_627) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_684) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_4_4) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_3) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_2) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_1) begin
          astInteract_4 <= 1'h0;
        end else if (kill_4_0) begin
          astInteract_4 <= 1'h0;
        end else if (_T_511) begin
          astInteract_4 <= _GEN_335;
        end else begin
          astInteract_4 <= _GEN_16;
        end
      end else begin
        astInteract_4 <= _GEN_16;
      end
    end else if (_T_862) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_886) begin
      astInteract_4 <= _GEN_16;
    end else if (_T_977) begin
      if (die_4) begin
        if (_T_1136) begin
          astInteract_4 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_4 <= 1'h0;
        end else begin
          astInteract_4 <= _GEN_16;
        end
      end else if (_T_1085) begin
        astInteract_4 <= 1'h0;
      end else begin
        astInteract_4 <= _GEN_16;
      end
    end else begin
      astInteract_4 <= _GEN_16;
    end
    if (reset) begin
      astInteract_5 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_5 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_505) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_570) begin
      if (kill_5_4) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_3) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_2) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_1) begin
        astInteract_5 <= 1'h0;
      end else if (kill_5_0) begin
        astInteract_5 <= 1'h0;
      end else if (_T_511) begin
        astInteract_5 <= _GEN_385;
      end else begin
        astInteract_5 <= _GEN_18;
      end
    end else if (_T_627) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_684) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_5_4) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_3) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_2) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_1) begin
          astInteract_5 <= 1'h0;
        end else if (kill_5_0) begin
          astInteract_5 <= 1'h0;
        end else if (_T_511) begin
          astInteract_5 <= _GEN_385;
        end else begin
          astInteract_5 <= _GEN_18;
        end
      end else begin
        astInteract_5 <= _GEN_18;
      end
    end else if (_T_862) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_886) begin
      astInteract_5 <= _GEN_18;
    end else if (_T_977) begin
      if (die_5) begin
        if (_T_1136) begin
          astInteract_5 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_5 <= 1'h0;
        end else begin
          astInteract_5 <= _GEN_18;
        end
      end else if (_T_1085) begin
        astInteract_5 <= 1'h0;
      end else begin
        astInteract_5 <= _GEN_18;
      end
    end else begin
      astInteract_5 <= _GEN_18;
    end
    if (reset) begin
      astInteract_6 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_6 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_505) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_570) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_627) begin
      if (kill_6_4) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_3) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_2) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_1) begin
        astInteract_6 <= 1'h0;
      end else if (kill_6_0) begin
        astInteract_6 <= 1'h0;
      end else if (_T_511) begin
        astInteract_6 <= _GEN_435;
      end else begin
        astInteract_6 <= _GEN_20;
      end
    end else if (_T_684) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_705) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_862) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_886) begin
      astInteract_6 <= _GEN_20;
    end else if (_T_977) begin
      if (die_6) begin
        if (_T_1136) begin
          astInteract_6 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_6 <= 1'h0;
        end else begin
          astInteract_6 <= _GEN_20;
        end
      end else if (_T_1085) begin
        astInteract_6 <= 1'h0;
      end else begin
        astInteract_6 <= _GEN_20;
      end
    end else begin
      astInteract_6 <= _GEN_20;
    end
    if (reset) begin
      astInteract_7 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_7 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_505) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_570) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_627) begin
      if (kill_7_4) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_3) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_2) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_1) begin
        astInteract_7 <= 1'h0;
      end else if (kill_7_0) begin
        astInteract_7 <= 1'h0;
      end else if (_T_511) begin
        astInteract_7 <= _GEN_485;
      end else begin
        astInteract_7 <= _GEN_22;
      end
    end else if (_T_684) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_705) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_862) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_886) begin
      astInteract_7 <= _GEN_22;
    end else if (_T_977) begin
      if (die_7) begin
        if (_T_1136) begin
          astInteract_7 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_7 <= 1'h0;
        end else begin
          astInteract_7 <= _GEN_22;
        end
      end else if (_T_1085) begin
        astInteract_7 <= 1'h0;
      end else begin
        astInteract_7 <= _GEN_22;
      end
    end else begin
      astInteract_7 <= _GEN_22;
    end
    if (reset) begin
      astInteract_8 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_8 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_505) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_570) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_627) begin
      if (kill_8_4) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_3) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_2) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_1) begin
        astInteract_8 <= 1'h0;
      end else if (kill_8_0) begin
        astInteract_8 <= 1'h0;
      end else if (_T_511) begin
        astInteract_8 <= _GEN_535;
      end else begin
        astInteract_8 <= _GEN_24;
      end
    end else if (_T_684) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_705) begin
      astInteract_8 <= 1'h0;
    end else if (_T_862) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_886) begin
      astInteract_8 <= _GEN_24;
    end else if (_T_977) begin
      if (die_8) begin
        if (_T_1136) begin
          astInteract_8 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_8 <= 1'h0;
        end else begin
          astInteract_8 <= _GEN_24;
        end
      end else if (_T_1085) begin
        astInteract_8 <= 1'h0;
      end else begin
        astInteract_8 <= _GEN_24;
      end
    end else begin
      astInteract_8 <= _GEN_24;
    end
    if (reset) begin
      astInteract_9 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_9 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_505) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_570) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_627) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_684) begin
      if (kill_9_3) begin
        astInteract_9 <= 1'h0;
      end else if (_T_688) begin
        astInteract_9 <= _GEN_585;
      end else begin
        astInteract_9 <= _GEN_26;
      end
    end else if (_T_705) begin
      if (_T_706) begin
        if (kill_9_3) begin
          astInteract_9 <= 1'h0;
        end else if (_T_688) begin
          astInteract_9 <= _GEN_585;
        end else begin
          astInteract_9 <= _GEN_26;
        end
      end else begin
        astInteract_9 <= _GEN_26;
      end
    end else if (_T_862) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_886) begin
      astInteract_9 <= _GEN_26;
    end else if (_T_977) begin
      if (die_9) begin
        if (_T_1136) begin
          astInteract_9 <= 1'h0;
        end else if (_T_1085) begin
          astInteract_9 <= 1'h0;
        end else begin
          astInteract_9 <= _GEN_26;
        end
      end else if (_T_1085) begin
        astInteract_9 <= 1'h0;
      end else begin
        astInteract_9 <= _GEN_26;
      end
    end else begin
      astInteract_9 <= _GEN_26;
    end
    if (reset) begin
      astInteract_10 <= 1'h0;
    end else if (_T_341) begin
      if (_T_340) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_342) begin
      if (_T_340) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_404) begin
      if (_T_340) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_451) begin
      if (_T_340) begin
        astInteract_10 <= 1'h0;
      end
    end else if (_T_486) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_505) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_570) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_627) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_684) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_705) begin
      if (_T_500) begin
        astInteract_10 <= 1'h0;
      end else if (_T_830) begin
        astInteract_10 <= _GEN_826;
      end else begin
        astInteract_10 <= _GEN_28;
      end
    end else if (_T_862) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_886) begin
      astInteract_10 <= _GEN_28;
    end else if (_T_977) begin
      if (die_10) begin
        if (_T_1136) begin
          astInteract_10 <= 1'h0;
        end else begin
          astInteract_10 <= _GEN_28;
        end
      end else begin
        astInteract_10 <= _GEN_28;
      end
    end else begin
      astInteract_10 <= _GEN_28;
    end
    shipInteract <= reset | _GEN_4255;
    if (reset) begin
      die_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_0 <= _T_1123;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_1 <= _T_1140;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_2 <= _T_1157;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_3 <= _T_1174;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_4 <= _T_1191;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_5 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_5 <= _T_1208;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_6 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_6 <= _T_1225;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_7 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_7 <= _T_1242;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_8 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_8 <= _T_1259;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_9 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_9 <= _T_1276;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      die_10 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              die_10 <= _T_1293;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_0_0 <= _T_1125;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_0_1 <= _T_1127;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_0_2 <= _T_1129;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_0_3 <= _T_1131;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_0_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_0_4 <= _T_1133;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_1_0 <= _T_1142;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_1_1 <= _T_1144;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_1_2 <= _T_1146;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_1_3 <= _T_1148;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_1_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_1_4 <= _T_1150;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_2_0 <= _T_1159;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_2_1 <= _T_1161;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_2_2 <= _T_1163;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_2_3 <= _T_1165;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_2_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_2_4 <= _T_1167;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_3_0 <= _T_1176;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_3_1 <= _T_1178;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_3_2 <= _T_1180;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_3_3 <= _T_1182;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_3_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_3_4 <= _T_1184;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_4_0 <= _T_1193;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_4_1 <= _T_1195;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_4_2 <= _T_1197;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_4_3 <= _T_1199;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_4_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_4_4 <= _T_1201;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_5_0 <= _T_1210;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_5_1 <= _T_1212;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_5_2 <= _T_1214;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_5_3 <= _T_1216;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_5_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_5_4 <= _T_1218;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_6_0 <= _T_1227;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_6_1 <= _T_1229;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_6_2 <= _T_1231;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_6_3 <= _T_1233;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_6_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_6_4 <= _T_1235;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_7_0 <= _T_1244;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_7_1 <= _T_1246;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_7_2 <= _T_1248;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_7_3 <= _T_1250;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_7_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_7_4 <= _T_1252;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_8_0 <= _T_1261;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_8_1 <= _T_1263;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_8_2 <= _T_1265;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_8_3 <= _T_1267;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_8_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_8_4 <= _T_1269;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_9_0 <= _T_1278;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_9_1 <= _T_1280;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_9_2 <= _T_1282;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_9_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_9_3 <= _T_1284;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_0 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_10_0 <= _T_1295;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_1 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_10_1 <= _T_1297;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_2 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_10_2 <= _T_1299;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_3 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_10_3 <= _T_1301;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      kill_10_4 <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              kill_10_4 <= _T_1303;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      hp <= 4'h3;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (io_sw_0) begin
                                hp <= 4'h3;
                              end else if (die_10) begin
                                if (_T_1136) begin
                                  hp <= _T_1138;
                                end else if (die_9) begin
                                  if (_T_1136) begin
                                    hp <= _T_1138;
                                  end else if (die_8) begin
                                    if (_T_1136) begin
                                      hp <= _T_1138;
                                    end else if (die_7) begin
                                      if (_T_1136) begin
                                        hp <= _T_1138;
                                      end else if (die_6) begin
                                        if (_T_1136) begin
                                          hp <= _T_1138;
                                        end else if (die_5) begin
                                          if (_T_1136) begin
                                            hp <= _T_1138;
                                          end else if (die_4) begin
                                            if (_T_1136) begin
                                              hp <= _T_1138;
                                            end else if (die_3) begin
                                              if (_T_1136) begin
                                                hp <= _T_1138;
                                              end else if (die_2) begin
                                                if (_T_1136) begin
                                                  hp <= _T_1138;
                                                end else if (die_1) begin
                                                  if (_T_1136) begin
                                                    hp <= _T_1138;
                                                  end else if (die_0) begin
                                                    if (_T_1136) begin
                                                      hp <= _T_1138;
                                                    end else if (_T_1088) begin
                                                      if (_T_1099) begin
                                                        hp <= 4'h3;
                                                      end
                                                    end
                                                  end else if (_T_1088) begin
                                                    if (_T_1099) begin
                                                      hp <= 4'h3;
                                                    end
                                                  end
                                                end else if (die_0) begin
                                                  if (_T_1136) begin
                                                    hp <= _T_1138;
                                                  end else if (_T_1088) begin
                                                    if (_T_1099) begin
                                                      hp <= 4'h3;
                                                    end
                                                  end
                                                end else if (_T_1088) begin
                                                  if (_T_1099) begin
                                                    hp <= 4'h3;
                                                  end
                                                end
                                              end else if (die_1) begin
                                                if (_T_1136) begin
                                                  hp <= _T_1138;
                                                end else if (die_0) begin
                                                  if (_T_1136) begin
                                                    hp <= _T_1138;
                                                  end else begin
                                                    hp <= _GEN_1169;
                                                  end
                                                end else begin
                                                  hp <= _GEN_1169;
                                                end
                                              end else if (die_0) begin
                                                if (_T_1136) begin
                                                  hp <= _T_1138;
                                                end else begin
                                                  hp <= _GEN_1169;
                                                end
                                              end else begin
                                                hp <= _GEN_1169;
                                              end
                                            end else if (die_2) begin
                                              if (_T_1136) begin
                                                hp <= _T_1138;
                                              end else if (die_1) begin
                                                if (_T_1136) begin
                                                  hp <= _T_1138;
                                                end else begin
                                                  hp <= _GEN_1184;
                                                end
                                              end else begin
                                                hp <= _GEN_1184;
                                              end
                                            end else if (die_1) begin
                                              if (_T_1136) begin
                                                hp <= _T_1138;
                                              end else begin
                                                hp <= _GEN_1184;
                                              end
                                            end else begin
                                              hp <= _GEN_1184;
                                            end
                                          end else if (die_3) begin
                                            if (_T_1136) begin
                                              hp <= _T_1138;
                                            end else if (die_2) begin
                                              if (_T_1136) begin
                                                hp <= _T_1138;
                                              end else begin
                                                hp <= _GEN_1194;
                                              end
                                            end else begin
                                              hp <= _GEN_1194;
                                            end
                                          end else if (die_2) begin
                                            if (_T_1136) begin
                                              hp <= _T_1138;
                                            end else begin
                                              hp <= _GEN_1194;
                                            end
                                          end else begin
                                            hp <= _GEN_1194;
                                          end
                                        end else if (die_4) begin
                                          if (_T_1136) begin
                                            hp <= _T_1138;
                                          end else if (die_3) begin
                                            if (_T_1136) begin
                                              hp <= _T_1138;
                                            end else begin
                                              hp <= _GEN_1204;
                                            end
                                          end else begin
                                            hp <= _GEN_1204;
                                          end
                                        end else if (die_3) begin
                                          if (_T_1136) begin
                                            hp <= _T_1138;
                                          end else begin
                                            hp <= _GEN_1204;
                                          end
                                        end else begin
                                          hp <= _GEN_1204;
                                        end
                                      end else if (die_5) begin
                                        if (_T_1136) begin
                                          hp <= _T_1138;
                                        end else if (die_4) begin
                                          if (_T_1136) begin
                                            hp <= _T_1138;
                                          end else begin
                                            hp <= _GEN_1214;
                                          end
                                        end else begin
                                          hp <= _GEN_1214;
                                        end
                                      end else if (die_4) begin
                                        if (_T_1136) begin
                                          hp <= _T_1138;
                                        end else begin
                                          hp <= _GEN_1214;
                                        end
                                      end else begin
                                        hp <= _GEN_1214;
                                      end
                                    end else if (die_6) begin
                                      if (_T_1136) begin
                                        hp <= _T_1138;
                                      end else if (die_5) begin
                                        if (_T_1136) begin
                                          hp <= _T_1138;
                                        end else begin
                                          hp <= _GEN_1224;
                                        end
                                      end else begin
                                        hp <= _GEN_1224;
                                      end
                                    end else if (die_5) begin
                                      if (_T_1136) begin
                                        hp <= _T_1138;
                                      end else begin
                                        hp <= _GEN_1224;
                                      end
                                    end else begin
                                      hp <= _GEN_1224;
                                    end
                                  end else if (die_7) begin
                                    if (_T_1136) begin
                                      hp <= _T_1138;
                                    end else if (die_6) begin
                                      if (_T_1136) begin
                                        hp <= _T_1138;
                                      end else begin
                                        hp <= _GEN_1234;
                                      end
                                    end else begin
                                      hp <= _GEN_1234;
                                    end
                                  end else if (die_6) begin
                                    if (_T_1136) begin
                                      hp <= _T_1138;
                                    end else begin
                                      hp <= _GEN_1234;
                                    end
                                  end else begin
                                    hp <= _GEN_1234;
                                  end
                                end else if (die_8) begin
                                  if (_T_1136) begin
                                    hp <= _T_1138;
                                  end else if (die_7) begin
                                    if (_T_1136) begin
                                      hp <= _T_1138;
                                    end else begin
                                      hp <= _GEN_1244;
                                    end
                                  end else begin
                                    hp <= _GEN_1244;
                                  end
                                end else if (die_7) begin
                                  if (_T_1136) begin
                                    hp <= _T_1138;
                                  end else begin
                                    hp <= _GEN_1244;
                                  end
                                end else begin
                                  hp <= _GEN_1244;
                                end
                              end else if (die_9) begin
                                if (_T_1136) begin
                                  hp <= _T_1138;
                                end else if (die_8) begin
                                  if (_T_1136) begin
                                    hp <= _T_1138;
                                  end else begin
                                    hp <= _GEN_1254;
                                  end
                                end else begin
                                  hp <= _GEN_1254;
                                end
                              end else if (die_8) begin
                                if (_T_1136) begin
                                  hp <= _T_1138;
                                end else begin
                                  hp <= _GEN_1254;
                                end
                              end else begin
                                hp <= _GEN_1254;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      planetHp <= 5'ha;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (_T_705) begin
                        if (kill_10_4) begin
                          if (_T_688) begin
                            planetHp <= _T_848;
                          end else if (kill_10_3) begin
                            if (_T_688) begin
                              planetHp <= _T_848;
                            end else if (kill_10_2) begin
                              if (_T_688) begin
                                planetHp <= _T_848;
                              end else if (kill_10_1) begin
                                if (_T_688) begin
                                  planetHp <= _T_848;
                                end else if (kill_10_0) begin
                                  if (_T_688) begin
                                    planetHp <= _T_848;
                                  end
                                end
                              end else if (kill_10_0) begin
                                if (_T_688) begin
                                  planetHp <= _T_848;
                                end
                              end
                            end else if (kill_10_1) begin
                              if (_T_688) begin
                                planetHp <= _T_848;
                              end else if (kill_10_0) begin
                                if (_T_688) begin
                                  planetHp <= _T_848;
                                end
                              end
                            end else if (kill_10_0) begin
                              if (_T_688) begin
                                planetHp <= _T_848;
                              end
                            end
                          end else if (kill_10_2) begin
                            if (_T_688) begin
                              planetHp <= _T_848;
                            end else if (kill_10_1) begin
                              if (_T_688) begin
                                planetHp <= _T_848;
                              end else begin
                                planetHp <= _GEN_835;
                              end
                            end else begin
                              planetHp <= _GEN_835;
                            end
                          end else if (kill_10_1) begin
                            if (_T_688) begin
                              planetHp <= _T_848;
                            end else begin
                              planetHp <= _GEN_835;
                            end
                          end else begin
                            planetHp <= _GEN_835;
                          end
                        end else if (kill_10_3) begin
                          if (_T_688) begin
                            planetHp <= _T_848;
                          end else if (kill_10_2) begin
                            if (_T_688) begin
                              planetHp <= _T_848;
                            end else begin
                              planetHp <= _GEN_840;
                            end
                          end else begin
                            planetHp <= _GEN_840;
                          end
                        end else if (kill_10_2) begin
                          if (_T_688) begin
                            planetHp <= _T_848;
                          end else begin
                            planetHp <= _GEN_840;
                          end
                        end else begin
                          planetHp <= _GEN_840;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      spwnProt <= 6'sh0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1314) begin
                                spwnProt <= 6'sh0;
                              end else if (_T_1310) begin
                                spwnProt <= _T_1313;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    show <= reset | _GEN_4246;
    if (reset) begin
      blink <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              blink <= _T_1116;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      secCnt <= 8'sh0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1088) begin
                                if (_T_1099) begin
                                  secCnt <= 8'sh0;
                                end else if (_T_1104) begin
                                  secCnt <= 8'shf;
                                end else begin
                                  secCnt <= _T_1091;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      level <= 3'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1088) begin
                                if (_T_1099) begin
                                  level <= _T_1101;
                                end else if (_T_500) begin
                                  level <= 3'h5;
                                end
                              end else if (_T_500) begin
                                level <= 3'h5;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      start <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              start <= _GEN_1294;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      levelCng <= 1'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (_T_404) begin
          if (_T_405) begin
            levelCng <= 1'h0;
          end
        end else if (!(_T_451)) begin
          if (!(_T_486)) begin
            if (!(_T_505)) begin
              if (!(_T_570)) begin
                if (!(_T_627)) begin
                  if (!(_T_684)) begin
                    if (!(_T_705)) begin
                      if (!(_T_862)) begin
                        if (!(_T_886)) begin
                          if (_T_977) begin
                            if (_T_1088) begin
                              levelCng <= _GEN_1167;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cngCnt <= 4'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1118) begin
                                if (_T_1121) begin
                                  cngCnt <= 4'h0;
                                end else begin
                                  cngCnt <= _T_1120;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cnt <= 10'sh0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1087) begin
                                cnt <= 10'sh0;
                              end else begin
                                cnt <= _T_1108;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      count1 <= 7'h0;
    end else if (!(_T_341)) begin
      if (_T_342) begin
        if (_T_395) begin
          if (levelCng) begin
            count1 <= _T_403;
          end
        end
      end else if (_T_404) begin
        if (_T_405) begin
          count1 <= 7'h0;
        end
      end else if (_T_451) begin
        if (_T_406) begin
          if (_T_407) begin
            count1 <= _T_403;
          end
        end
      end
    end
    if (reset) begin
      count3 <= 7'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (_T_404) begin
          if (_T_437) begin
            if (_T_408) begin
              count3 <= _T_420;
            end else begin
              count3 <= 7'h0;
            end
          end else if (_T_423) begin
            if (_T_408) begin
              count3 <= _T_420;
            end else begin
              count3 <= 7'h0;
            end
          end else if (_T_406) begin
            if (_T_407) begin
              if (_T_408) begin
                count3 <= _T_420;
              end else begin
                count3 <= 7'h0;
              end
            end
          end
        end else if (_T_451) begin
          if (_T_437) begin
            if (_T_408) begin
              count3 <= _T_420;
            end else begin
              count3 <= 7'h0;
            end
          end else if (_T_423) begin
            count3 <= _GEN_40;
          end
        end else if (_T_486) begin
          if (_T_408) begin
            count3 <= _T_420;
          end else if (!(_T_500)) begin
            count3 <= 7'h0;
          end
        end
      end
    end
    if (reset) begin
      count4 <= 8'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (_T_451) begin
            if (_T_423) begin
              if (_T_408) begin
                if (_T_406) begin
                  if (_T_407) begin
                    count4 <= 8'h0;
                  end
                end
              end else begin
                count4 <= 8'h1;
              end
            end else if (_T_406) begin
              if (_T_407) begin
                count4 <= 8'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      count5 <= 8'h0;
    end else if (!(_T_341)) begin
      if (!(_T_342)) begin
        if (!(_T_404)) begin
          if (!(_T_451)) begin
            if (!(_T_486)) begin
              if (!(_T_505)) begin
                if (!(_T_570)) begin
                  if (!(_T_627)) begin
                    if (!(_T_684)) begin
                      if (!(_T_705)) begin
                        if (!(_T_862)) begin
                          if (!(_T_886)) begin
                            if (_T_977) begin
                              if (_T_1026) begin
                                count5 <= 8'h1;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    _T_912 <= Xstart_0;
    _T_917 <= Ystart_0;
    _T_927 <= Xstart_0;
    _T_932 <= Ystart_0;
    _T_940 <= Xstart_0;
    _T_945 <= Ystart_0;
    _T_953 <= Xstart_0;
    _T_958 <= Ystart_0;
    _T_966 <= Xstart_0;
    _T_971 <= Ystart_0;
    if (reset) begin
      _T_978 <= 1'h0;
    end else begin
      _T_978 <= _GEN_1078;
    end
    if (reset) begin
      _T_979 <= 1'h0;
    end else begin
      _T_979 <= _GEN_1079;
    end
    if (reset) begin
      _T_980 <= 3'sh0;
    end else if (_T_983) begin
      _T_980 <= {{1{Randomizer_33_io_out[1]}},Randomizer_33_io_out};
    end
    if (reset) begin
      _T_981 <= 3'sh0;
    end else if (_T_984) begin
      _T_981 <= {{1{Randomizer_33_io_out[1]}},Randomizer_33_io_out};
    end
    if (reset) begin
      _T_982 <= 3'sh0;
    end else if (_T_985) begin
      _T_982 <= {{1{Randomizer_33_io_out[1]}},Randomizer_33_io_out};
    end
    if (reset) begin
      _T_1028 <= 1'h0;
    end else begin
      _T_1028 <= _GEN_1107;
    end
    if (reset) begin
      _T_1029 <= 1'h0;
    end else begin
      _T_1029 <= _GEN_1108;
    end
    if (reset) begin
      _T_1030 <= 3'sh0;
    end else if (_T_1033) begin
      _T_1030 <= {{1{Randomizer_40_io_out[1]}},Randomizer_40_io_out};
    end
    if (reset) begin
      _T_1031 <= 3'sh0;
    end else if (_T_1034) begin
      _T_1031 <= {{1{Randomizer_40_io_out[1]}},Randomizer_40_io_out};
    end
    if (reset) begin
      _T_1032 <= 3'sh0;
    end else if (_T_1035) begin
      _T_1032 <= {{1{Randomizer_40_io_out[1]}},Randomizer_40_io_out};
    end
  end
endmodule
module GameTop(
  input        clock,
  input        reset,
  input        io_btnC,
  input        io_btnU,
  input        io_btnL,
  input        io_btnR,
  input        io_btnD,
  output [3:0] io_vgaRed,
  output [3:0] io_vgaBlue,
  output [3:0] io_vgaGreen,
  output       io_Hsync,
  output       io_Vsync,
  input        io_sw_0,
  input        io_sw_1,
  input        io_sw_2,
  input        io_sw_7,
  output       io_soundOutput_0,
  output       io_missingFrameError,
  output       io_backBufferWriteError,
  output       io_viewBoxOutOfRangeError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire  graphicEngineVGA_clock; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_reset; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_0; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_1; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_2; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_3; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_4; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_5; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_6; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_7; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_8; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_9; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_10; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_11; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_12; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_13; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_14; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_15; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_16; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_17; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_18; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_19; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_20; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_21; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_22; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_23; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_24; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_25; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_26; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_27; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_28; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_29; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_30; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_31; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_32; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_33; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_41; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_42; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_43; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_44; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_45; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_46; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_47; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_48; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_49; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_50; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_51; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_122; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_123; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_124; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_125; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_126; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_spriteXPosition_127; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_0; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_1; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_2; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_3; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_4; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_5; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_6; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_7; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_8; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_9; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_10; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_11; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_12; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_13; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_14; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_15; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_16; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_17; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_18; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_19; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_20; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_21; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_22; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_23; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_24; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_25; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_26; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_27; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_28; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_29; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_30; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_31; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_32; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_33; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_41; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_42; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_43; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_122; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_123; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_124; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_125; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_126; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_spriteYPosition_127; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_0; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_1; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_2; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_3; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_4; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_5; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_6; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_7; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_8; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_9; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_10; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_11; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_12; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_13; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_14; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_15; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_16; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_17; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_18; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_19; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_20; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_21; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_22; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_23; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_24; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_25; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_26; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_27; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_28; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_29; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_30; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_31; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_32; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_33; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_41; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_42; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_43; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_44; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_45; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_46; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_47; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_48; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_49; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_50; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_51; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_55; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_56; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_57; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_61; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_62; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_63; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_64; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_65; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_66; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_70; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_71; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteVisible_72; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_122; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_123; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_124; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_125; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_126; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_spriteFlipVertical_127; // @[GameTop.scala 46:32]
  wire [9:0] graphicEngineVGA_io_viewBoxX_0; // @[GameTop.scala 46:32]
  wire [4:0] graphicEngineVGA_io_backBufferWriteData; // @[GameTop.scala 46:32]
  wire [10:0] graphicEngineVGA_io_backBufferWriteAddress; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_backBufferWriteEnable; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_newFrame; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_frameUpdateDone; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_missingFrameError; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_backBufferWriteError; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_viewBoxOutOfRangeError; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaRed; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaBlue; // @[GameTop.scala 46:32]
  wire [3:0] graphicEngineVGA_io_vgaGreen; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Hsync; // @[GameTop.scala 46:32]
  wire  graphicEngineVGA_io_Vsync; // @[GameTop.scala 46:32]
  wire  soundEngine_clock; // @[GameTop.scala 48:27]
  wire  soundEngine_reset; // @[GameTop.scala 48:27]
  wire  soundEngine_io_output_0; // @[GameTop.scala 48:27]
  wire [3:0] soundEngine_io_input; // @[GameTop.scala 48:27]
  wire  gameLogic_clock; // @[GameTop.scala 52:25]
  wire  gameLogic_reset; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnC; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnU; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnL; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnR; // @[GameTop.scala 52:25]
  wire  gameLogic_io_btnD; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_0; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_1; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_2; // @[GameTop.scala 52:25]
  wire  gameLogic_io_sw_7; // @[GameTop.scala 52:25]
  wire [3:0] gameLogic_io_songInput; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_0; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_1; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_2; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_3; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_4; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_5; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_6; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_7; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_8; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_9; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_10; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_11; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_12; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_13; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_14; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_15; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_16; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_17; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_18; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_19; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_20; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_21; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_22; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_23; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_24; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_25; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_26; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_27; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_28; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_29; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_30; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_31; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_32; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_33; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_41; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_42; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_43; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_44; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_45; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_46; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_47; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_48; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_49; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_50; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_51; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_122; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_123; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_124; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_125; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_126; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_spriteXPosition_127; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_0; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_1; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_2; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_3; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_4; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_5; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_6; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_7; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_8; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_9; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_10; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_11; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_12; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_13; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_14; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_15; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_16; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_17; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_18; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_19; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_20; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_21; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_22; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_23; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_24; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_25; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_26; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_27; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_28; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_29; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_30; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_31; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_32; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_33; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_41; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_42; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_43; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_122; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_123; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_124; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_125; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_126; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_spriteYPosition_127; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_0; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_1; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_2; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_3; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_4; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_5; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_6; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_7; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_8; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_9; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_10; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_11; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_12; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_13; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_14; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_15; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_16; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_17; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_18; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_19; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_20; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_21; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_22; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_23; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_24; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_25; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_26; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_27; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_28; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_29; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_30; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_31; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_32; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_33; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_41; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_42; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_43; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_44; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_45; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_46; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_47; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_48; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_49; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_50; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_51; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_55; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_56; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_57; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_61; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_62; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_63; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_64; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_65; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_66; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_70; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_71; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteVisible_72; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_122; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_123; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_124; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_125; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_126; // @[GameTop.scala 52:25]
  wire  gameLogic_io_spriteFlipVertical_127; // @[GameTop.scala 52:25]
  wire [9:0] gameLogic_io_viewBoxX_0; // @[GameTop.scala 52:25]
  wire [4:0] gameLogic_io_backBufferWriteData; // @[GameTop.scala 52:25]
  wire [10:0] gameLogic_io_backBufferWriteAddress; // @[GameTop.scala 52:25]
  wire  gameLogic_io_backBufferWriteEnable; // @[GameTop.scala 52:25]
  wire  gameLogic_io_newFrame; // @[GameTop.scala 52:25]
  wire  gameLogic_io_frameUpdateDone; // @[GameTop.scala 52:25]
  reg [20:0] debounceCounter; // @[GameTop.scala 72:32]
  wire  debounceSampleEn = debounceCounter == 21'h1e847f; // @[GameTop.scala 74:24]
  wire [20:0] _T_2 = debounceCounter + 21'h1; // @[GameTop.scala 78:40]
  reg [21:0] resetReleaseCounter; // @[GameTop.scala 85:36]
  wire  _T_3 = resetReleaseCounter == 22'h3d08ff; // @[GameTop.scala 87:28]
  wire [21:0] _T_5 = resetReleaseCounter + 22'h1; // @[GameTop.scala 91:48]
  reg  _T_7_0; // @[GameUtilities.scala 39:28]
  reg  _T_7_1; // @[GameUtilities.scala 39:28]
  reg  _T_7_2; // @[GameUtilities.scala 39:28]
  reg  btnCState; // @[Reg.scala 27:20]
  reg  _T_9_0; // @[GameUtilities.scala 39:28]
  reg  _T_9_1; // @[GameUtilities.scala 39:28]
  reg  _T_9_2; // @[GameUtilities.scala 39:28]
  reg  btnUState; // @[Reg.scala 27:20]
  reg  _T_11_0; // @[GameUtilities.scala 39:28]
  reg  _T_11_1; // @[GameUtilities.scala 39:28]
  reg  _T_11_2; // @[GameUtilities.scala 39:28]
  reg  btnLState; // @[Reg.scala 27:20]
  reg  _T_13_0; // @[GameUtilities.scala 39:28]
  reg  _T_13_1; // @[GameUtilities.scala 39:28]
  reg  _T_13_2; // @[GameUtilities.scala 39:28]
  reg  btnRState; // @[Reg.scala 27:20]
  reg  _T_15_0; // @[GameUtilities.scala 39:28]
  reg  _T_15_1; // @[GameUtilities.scala 39:28]
  reg  _T_15_2; // @[GameUtilities.scala 39:28]
  reg  btnDState; // @[Reg.scala 27:20]
  reg  _T_17_0; // @[GameUtilities.scala 39:28]
  reg  _T_17_1; // @[GameUtilities.scala 39:28]
  reg  _T_17_2; // @[GameUtilities.scala 39:28]
  reg  _T_18; // @[Reg.scala 27:20]
  reg  _T_20_0; // @[GameUtilities.scala 39:28]
  reg  _T_20_1; // @[GameUtilities.scala 39:28]
  reg  _T_20_2; // @[GameUtilities.scala 39:28]
  reg  _T_21; // @[Reg.scala 27:20]
  reg  _T_23_0; // @[GameUtilities.scala 39:28]
  reg  _T_23_1; // @[GameUtilities.scala 39:28]
  reg  _T_23_2; // @[GameUtilities.scala 39:28]
  reg  _T_24; // @[Reg.scala 27:20]
  reg  _T_38_0; // @[GameUtilities.scala 39:28]
  reg  _T_38_1; // @[GameUtilities.scala 39:28]
  reg  _T_38_2; // @[GameUtilities.scala 39:28]
  reg  _T_39; // @[Reg.scala 27:20]
  GraphicEngineVGA graphicEngineVGA ( // @[GameTop.scala 46:32]
    .clock(graphicEngineVGA_clock),
    .reset(graphicEngineVGA_reset),
    .io_spriteXPosition_0(graphicEngineVGA_io_spriteXPosition_0),
    .io_spriteXPosition_1(graphicEngineVGA_io_spriteXPosition_1),
    .io_spriteXPosition_2(graphicEngineVGA_io_spriteXPosition_2),
    .io_spriteXPosition_3(graphicEngineVGA_io_spriteXPosition_3),
    .io_spriteXPosition_4(graphicEngineVGA_io_spriteXPosition_4),
    .io_spriteXPosition_5(graphicEngineVGA_io_spriteXPosition_5),
    .io_spriteXPosition_6(graphicEngineVGA_io_spriteXPosition_6),
    .io_spriteXPosition_7(graphicEngineVGA_io_spriteXPosition_7),
    .io_spriteXPosition_8(graphicEngineVGA_io_spriteXPosition_8),
    .io_spriteXPosition_9(graphicEngineVGA_io_spriteXPosition_9),
    .io_spriteXPosition_10(graphicEngineVGA_io_spriteXPosition_10),
    .io_spriteXPosition_11(graphicEngineVGA_io_spriteXPosition_11),
    .io_spriteXPosition_12(graphicEngineVGA_io_spriteXPosition_12),
    .io_spriteXPosition_13(graphicEngineVGA_io_spriteXPosition_13),
    .io_spriteXPosition_14(graphicEngineVGA_io_spriteXPosition_14),
    .io_spriteXPosition_15(graphicEngineVGA_io_spriteXPosition_15),
    .io_spriteXPosition_16(graphicEngineVGA_io_spriteXPosition_16),
    .io_spriteXPosition_17(graphicEngineVGA_io_spriteXPosition_17),
    .io_spriteXPosition_18(graphicEngineVGA_io_spriteXPosition_18),
    .io_spriteXPosition_19(graphicEngineVGA_io_spriteXPosition_19),
    .io_spriteXPosition_20(graphicEngineVGA_io_spriteXPosition_20),
    .io_spriteXPosition_21(graphicEngineVGA_io_spriteXPosition_21),
    .io_spriteXPosition_22(graphicEngineVGA_io_spriteXPosition_22),
    .io_spriteXPosition_23(graphicEngineVGA_io_spriteXPosition_23),
    .io_spriteXPosition_24(graphicEngineVGA_io_spriteXPosition_24),
    .io_spriteXPosition_25(graphicEngineVGA_io_spriteXPosition_25),
    .io_spriteXPosition_26(graphicEngineVGA_io_spriteXPosition_26),
    .io_spriteXPosition_27(graphicEngineVGA_io_spriteXPosition_27),
    .io_spriteXPosition_28(graphicEngineVGA_io_spriteXPosition_28),
    .io_spriteXPosition_29(graphicEngineVGA_io_spriteXPosition_29),
    .io_spriteXPosition_30(graphicEngineVGA_io_spriteXPosition_30),
    .io_spriteXPosition_31(graphicEngineVGA_io_spriteXPosition_31),
    .io_spriteXPosition_32(graphicEngineVGA_io_spriteXPosition_32),
    .io_spriteXPosition_33(graphicEngineVGA_io_spriteXPosition_33),
    .io_spriteXPosition_41(graphicEngineVGA_io_spriteXPosition_41),
    .io_spriteXPosition_42(graphicEngineVGA_io_spriteXPosition_42),
    .io_spriteXPosition_43(graphicEngineVGA_io_spriteXPosition_43),
    .io_spriteXPosition_44(graphicEngineVGA_io_spriteXPosition_44),
    .io_spriteXPosition_45(graphicEngineVGA_io_spriteXPosition_45),
    .io_spriteXPosition_46(graphicEngineVGA_io_spriteXPosition_46),
    .io_spriteXPosition_47(graphicEngineVGA_io_spriteXPosition_47),
    .io_spriteXPosition_48(graphicEngineVGA_io_spriteXPosition_48),
    .io_spriteXPosition_49(graphicEngineVGA_io_spriteXPosition_49),
    .io_spriteXPosition_50(graphicEngineVGA_io_spriteXPosition_50),
    .io_spriteXPosition_51(graphicEngineVGA_io_spriteXPosition_51),
    .io_spriteXPosition_122(graphicEngineVGA_io_spriteXPosition_122),
    .io_spriteXPosition_123(graphicEngineVGA_io_spriteXPosition_123),
    .io_spriteXPosition_124(graphicEngineVGA_io_spriteXPosition_124),
    .io_spriteXPosition_125(graphicEngineVGA_io_spriteXPosition_125),
    .io_spriteXPosition_126(graphicEngineVGA_io_spriteXPosition_126),
    .io_spriteXPosition_127(graphicEngineVGA_io_spriteXPosition_127),
    .io_spriteYPosition_0(graphicEngineVGA_io_spriteYPosition_0),
    .io_spriteYPosition_1(graphicEngineVGA_io_spriteYPosition_1),
    .io_spriteYPosition_2(graphicEngineVGA_io_spriteYPosition_2),
    .io_spriteYPosition_3(graphicEngineVGA_io_spriteYPosition_3),
    .io_spriteYPosition_4(graphicEngineVGA_io_spriteYPosition_4),
    .io_spriteYPosition_5(graphicEngineVGA_io_spriteYPosition_5),
    .io_spriteYPosition_6(graphicEngineVGA_io_spriteYPosition_6),
    .io_spriteYPosition_7(graphicEngineVGA_io_spriteYPosition_7),
    .io_spriteYPosition_8(graphicEngineVGA_io_spriteYPosition_8),
    .io_spriteYPosition_9(graphicEngineVGA_io_spriteYPosition_9),
    .io_spriteYPosition_10(graphicEngineVGA_io_spriteYPosition_10),
    .io_spriteYPosition_11(graphicEngineVGA_io_spriteYPosition_11),
    .io_spriteYPosition_12(graphicEngineVGA_io_spriteYPosition_12),
    .io_spriteYPosition_13(graphicEngineVGA_io_spriteYPosition_13),
    .io_spriteYPosition_14(graphicEngineVGA_io_spriteYPosition_14),
    .io_spriteYPosition_15(graphicEngineVGA_io_spriteYPosition_15),
    .io_spriteYPosition_16(graphicEngineVGA_io_spriteYPosition_16),
    .io_spriteYPosition_17(graphicEngineVGA_io_spriteYPosition_17),
    .io_spriteYPosition_18(graphicEngineVGA_io_spriteYPosition_18),
    .io_spriteYPosition_19(graphicEngineVGA_io_spriteYPosition_19),
    .io_spriteYPosition_20(graphicEngineVGA_io_spriteYPosition_20),
    .io_spriteYPosition_21(graphicEngineVGA_io_spriteYPosition_21),
    .io_spriteYPosition_22(graphicEngineVGA_io_spriteYPosition_22),
    .io_spriteYPosition_23(graphicEngineVGA_io_spriteYPosition_23),
    .io_spriteYPosition_24(graphicEngineVGA_io_spriteYPosition_24),
    .io_spriteYPosition_25(graphicEngineVGA_io_spriteYPosition_25),
    .io_spriteYPosition_26(graphicEngineVGA_io_spriteYPosition_26),
    .io_spriteYPosition_27(graphicEngineVGA_io_spriteYPosition_27),
    .io_spriteYPosition_28(graphicEngineVGA_io_spriteYPosition_28),
    .io_spriteYPosition_29(graphicEngineVGA_io_spriteYPosition_29),
    .io_spriteYPosition_30(graphicEngineVGA_io_spriteYPosition_30),
    .io_spriteYPosition_31(graphicEngineVGA_io_spriteYPosition_31),
    .io_spriteYPosition_32(graphicEngineVGA_io_spriteYPosition_32),
    .io_spriteYPosition_33(graphicEngineVGA_io_spriteYPosition_33),
    .io_spriteYPosition_41(graphicEngineVGA_io_spriteYPosition_41),
    .io_spriteYPosition_42(graphicEngineVGA_io_spriteYPosition_42),
    .io_spriteYPosition_43(graphicEngineVGA_io_spriteYPosition_43),
    .io_spriteYPosition_122(graphicEngineVGA_io_spriteYPosition_122),
    .io_spriteYPosition_123(graphicEngineVGA_io_spriteYPosition_123),
    .io_spriteYPosition_124(graphicEngineVGA_io_spriteYPosition_124),
    .io_spriteYPosition_125(graphicEngineVGA_io_spriteYPosition_125),
    .io_spriteYPosition_126(graphicEngineVGA_io_spriteYPosition_126),
    .io_spriteYPosition_127(graphicEngineVGA_io_spriteYPosition_127),
    .io_spriteVisible_0(graphicEngineVGA_io_spriteVisible_0),
    .io_spriteVisible_1(graphicEngineVGA_io_spriteVisible_1),
    .io_spriteVisible_2(graphicEngineVGA_io_spriteVisible_2),
    .io_spriteVisible_3(graphicEngineVGA_io_spriteVisible_3),
    .io_spriteVisible_4(graphicEngineVGA_io_spriteVisible_4),
    .io_spriteVisible_5(graphicEngineVGA_io_spriteVisible_5),
    .io_spriteVisible_6(graphicEngineVGA_io_spriteVisible_6),
    .io_spriteVisible_7(graphicEngineVGA_io_spriteVisible_7),
    .io_spriteVisible_8(graphicEngineVGA_io_spriteVisible_8),
    .io_spriteVisible_9(graphicEngineVGA_io_spriteVisible_9),
    .io_spriteVisible_10(graphicEngineVGA_io_spriteVisible_10),
    .io_spriteVisible_11(graphicEngineVGA_io_spriteVisible_11),
    .io_spriteVisible_12(graphicEngineVGA_io_spriteVisible_12),
    .io_spriteVisible_13(graphicEngineVGA_io_spriteVisible_13),
    .io_spriteVisible_14(graphicEngineVGA_io_spriteVisible_14),
    .io_spriteVisible_15(graphicEngineVGA_io_spriteVisible_15),
    .io_spriteVisible_16(graphicEngineVGA_io_spriteVisible_16),
    .io_spriteVisible_17(graphicEngineVGA_io_spriteVisible_17),
    .io_spriteVisible_18(graphicEngineVGA_io_spriteVisible_18),
    .io_spriteVisible_19(graphicEngineVGA_io_spriteVisible_19),
    .io_spriteVisible_20(graphicEngineVGA_io_spriteVisible_20),
    .io_spriteVisible_21(graphicEngineVGA_io_spriteVisible_21),
    .io_spriteVisible_22(graphicEngineVGA_io_spriteVisible_22),
    .io_spriteVisible_23(graphicEngineVGA_io_spriteVisible_23),
    .io_spriteVisible_24(graphicEngineVGA_io_spriteVisible_24),
    .io_spriteVisible_25(graphicEngineVGA_io_spriteVisible_25),
    .io_spriteVisible_26(graphicEngineVGA_io_spriteVisible_26),
    .io_spriteVisible_27(graphicEngineVGA_io_spriteVisible_27),
    .io_spriteVisible_28(graphicEngineVGA_io_spriteVisible_28),
    .io_spriteVisible_29(graphicEngineVGA_io_spriteVisible_29),
    .io_spriteVisible_30(graphicEngineVGA_io_spriteVisible_30),
    .io_spriteVisible_31(graphicEngineVGA_io_spriteVisible_31),
    .io_spriteVisible_32(graphicEngineVGA_io_spriteVisible_32),
    .io_spriteVisible_33(graphicEngineVGA_io_spriteVisible_33),
    .io_spriteVisible_41(graphicEngineVGA_io_spriteVisible_41),
    .io_spriteVisible_42(graphicEngineVGA_io_spriteVisible_42),
    .io_spriteVisible_43(graphicEngineVGA_io_spriteVisible_43),
    .io_spriteVisible_44(graphicEngineVGA_io_spriteVisible_44),
    .io_spriteVisible_45(graphicEngineVGA_io_spriteVisible_45),
    .io_spriteVisible_46(graphicEngineVGA_io_spriteVisible_46),
    .io_spriteVisible_47(graphicEngineVGA_io_spriteVisible_47),
    .io_spriteVisible_48(graphicEngineVGA_io_spriteVisible_48),
    .io_spriteVisible_49(graphicEngineVGA_io_spriteVisible_49),
    .io_spriteVisible_50(graphicEngineVGA_io_spriteVisible_50),
    .io_spriteVisible_51(graphicEngineVGA_io_spriteVisible_51),
    .io_spriteVisible_55(graphicEngineVGA_io_spriteVisible_55),
    .io_spriteVisible_56(graphicEngineVGA_io_spriteVisible_56),
    .io_spriteVisible_57(graphicEngineVGA_io_spriteVisible_57),
    .io_spriteVisible_61(graphicEngineVGA_io_spriteVisible_61),
    .io_spriteVisible_62(graphicEngineVGA_io_spriteVisible_62),
    .io_spriteVisible_63(graphicEngineVGA_io_spriteVisible_63),
    .io_spriteVisible_64(graphicEngineVGA_io_spriteVisible_64),
    .io_spriteVisible_65(graphicEngineVGA_io_spriteVisible_65),
    .io_spriteVisible_66(graphicEngineVGA_io_spriteVisible_66),
    .io_spriteVisible_70(graphicEngineVGA_io_spriteVisible_70),
    .io_spriteVisible_71(graphicEngineVGA_io_spriteVisible_71),
    .io_spriteVisible_72(graphicEngineVGA_io_spriteVisible_72),
    .io_spriteFlipVertical_122(graphicEngineVGA_io_spriteFlipVertical_122),
    .io_spriteFlipVertical_123(graphicEngineVGA_io_spriteFlipVertical_123),
    .io_spriteFlipVertical_124(graphicEngineVGA_io_spriteFlipVertical_124),
    .io_spriteFlipVertical_125(graphicEngineVGA_io_spriteFlipVertical_125),
    .io_spriteFlipVertical_126(graphicEngineVGA_io_spriteFlipVertical_126),
    .io_spriteFlipVertical_127(graphicEngineVGA_io_spriteFlipVertical_127),
    .io_viewBoxX_0(graphicEngineVGA_io_viewBoxX_0),
    .io_backBufferWriteData(graphicEngineVGA_io_backBufferWriteData),
    .io_backBufferWriteAddress(graphicEngineVGA_io_backBufferWriteAddress),
    .io_backBufferWriteEnable(graphicEngineVGA_io_backBufferWriteEnable),
    .io_newFrame(graphicEngineVGA_io_newFrame),
    .io_frameUpdateDone(graphicEngineVGA_io_frameUpdateDone),
    .io_missingFrameError(graphicEngineVGA_io_missingFrameError),
    .io_backBufferWriteError(graphicEngineVGA_io_backBufferWriteError),
    .io_viewBoxOutOfRangeError(graphicEngineVGA_io_viewBoxOutOfRangeError),
    .io_vgaRed(graphicEngineVGA_io_vgaRed),
    .io_vgaBlue(graphicEngineVGA_io_vgaBlue),
    .io_vgaGreen(graphicEngineVGA_io_vgaGreen),
    .io_Hsync(graphicEngineVGA_io_Hsync),
    .io_Vsync(graphicEngineVGA_io_Vsync)
  );
  SoundEngine soundEngine ( // @[GameTop.scala 48:27]
    .clock(soundEngine_clock),
    .reset(soundEngine_reset),
    .io_output_0(soundEngine_io_output_0),
    .io_input(soundEngine_io_input)
  );
  GameLogic gameLogic ( // @[GameTop.scala 52:25]
    .clock(gameLogic_clock),
    .reset(gameLogic_reset),
    .io_btnC(gameLogic_io_btnC),
    .io_btnU(gameLogic_io_btnU),
    .io_btnL(gameLogic_io_btnL),
    .io_btnR(gameLogic_io_btnR),
    .io_btnD(gameLogic_io_btnD),
    .io_sw_0(gameLogic_io_sw_0),
    .io_sw_1(gameLogic_io_sw_1),
    .io_sw_2(gameLogic_io_sw_2),
    .io_sw_7(gameLogic_io_sw_7),
    .io_songInput(gameLogic_io_songInput),
    .io_spriteXPosition_0(gameLogic_io_spriteXPosition_0),
    .io_spriteXPosition_1(gameLogic_io_spriteXPosition_1),
    .io_spriteXPosition_2(gameLogic_io_spriteXPosition_2),
    .io_spriteXPosition_3(gameLogic_io_spriteXPosition_3),
    .io_spriteXPosition_4(gameLogic_io_spriteXPosition_4),
    .io_spriteXPosition_5(gameLogic_io_spriteXPosition_5),
    .io_spriteXPosition_6(gameLogic_io_spriteXPosition_6),
    .io_spriteXPosition_7(gameLogic_io_spriteXPosition_7),
    .io_spriteXPosition_8(gameLogic_io_spriteXPosition_8),
    .io_spriteXPosition_9(gameLogic_io_spriteXPosition_9),
    .io_spriteXPosition_10(gameLogic_io_spriteXPosition_10),
    .io_spriteXPosition_11(gameLogic_io_spriteXPosition_11),
    .io_spriteXPosition_12(gameLogic_io_spriteXPosition_12),
    .io_spriteXPosition_13(gameLogic_io_spriteXPosition_13),
    .io_spriteXPosition_14(gameLogic_io_spriteXPosition_14),
    .io_spriteXPosition_15(gameLogic_io_spriteXPosition_15),
    .io_spriteXPosition_16(gameLogic_io_spriteXPosition_16),
    .io_spriteXPosition_17(gameLogic_io_spriteXPosition_17),
    .io_spriteXPosition_18(gameLogic_io_spriteXPosition_18),
    .io_spriteXPosition_19(gameLogic_io_spriteXPosition_19),
    .io_spriteXPosition_20(gameLogic_io_spriteXPosition_20),
    .io_spriteXPosition_21(gameLogic_io_spriteXPosition_21),
    .io_spriteXPosition_22(gameLogic_io_spriteXPosition_22),
    .io_spriteXPosition_23(gameLogic_io_spriteXPosition_23),
    .io_spriteXPosition_24(gameLogic_io_spriteXPosition_24),
    .io_spriteXPosition_25(gameLogic_io_spriteXPosition_25),
    .io_spriteXPosition_26(gameLogic_io_spriteXPosition_26),
    .io_spriteXPosition_27(gameLogic_io_spriteXPosition_27),
    .io_spriteXPosition_28(gameLogic_io_spriteXPosition_28),
    .io_spriteXPosition_29(gameLogic_io_spriteXPosition_29),
    .io_spriteXPosition_30(gameLogic_io_spriteXPosition_30),
    .io_spriteXPosition_31(gameLogic_io_spriteXPosition_31),
    .io_spriteXPosition_32(gameLogic_io_spriteXPosition_32),
    .io_spriteXPosition_33(gameLogic_io_spriteXPosition_33),
    .io_spriteXPosition_41(gameLogic_io_spriteXPosition_41),
    .io_spriteXPosition_42(gameLogic_io_spriteXPosition_42),
    .io_spriteXPosition_43(gameLogic_io_spriteXPosition_43),
    .io_spriteXPosition_44(gameLogic_io_spriteXPosition_44),
    .io_spriteXPosition_45(gameLogic_io_spriteXPosition_45),
    .io_spriteXPosition_46(gameLogic_io_spriteXPosition_46),
    .io_spriteXPosition_47(gameLogic_io_spriteXPosition_47),
    .io_spriteXPosition_48(gameLogic_io_spriteXPosition_48),
    .io_spriteXPosition_49(gameLogic_io_spriteXPosition_49),
    .io_spriteXPosition_50(gameLogic_io_spriteXPosition_50),
    .io_spriteXPosition_51(gameLogic_io_spriteXPosition_51),
    .io_spriteXPosition_122(gameLogic_io_spriteXPosition_122),
    .io_spriteXPosition_123(gameLogic_io_spriteXPosition_123),
    .io_spriteXPosition_124(gameLogic_io_spriteXPosition_124),
    .io_spriteXPosition_125(gameLogic_io_spriteXPosition_125),
    .io_spriteXPosition_126(gameLogic_io_spriteXPosition_126),
    .io_spriteXPosition_127(gameLogic_io_spriteXPosition_127),
    .io_spriteYPosition_0(gameLogic_io_spriteYPosition_0),
    .io_spriteYPosition_1(gameLogic_io_spriteYPosition_1),
    .io_spriteYPosition_2(gameLogic_io_spriteYPosition_2),
    .io_spriteYPosition_3(gameLogic_io_spriteYPosition_3),
    .io_spriteYPosition_4(gameLogic_io_spriteYPosition_4),
    .io_spriteYPosition_5(gameLogic_io_spriteYPosition_5),
    .io_spriteYPosition_6(gameLogic_io_spriteYPosition_6),
    .io_spriteYPosition_7(gameLogic_io_spriteYPosition_7),
    .io_spriteYPosition_8(gameLogic_io_spriteYPosition_8),
    .io_spriteYPosition_9(gameLogic_io_spriteYPosition_9),
    .io_spriteYPosition_10(gameLogic_io_spriteYPosition_10),
    .io_spriteYPosition_11(gameLogic_io_spriteYPosition_11),
    .io_spriteYPosition_12(gameLogic_io_spriteYPosition_12),
    .io_spriteYPosition_13(gameLogic_io_spriteYPosition_13),
    .io_spriteYPosition_14(gameLogic_io_spriteYPosition_14),
    .io_spriteYPosition_15(gameLogic_io_spriteYPosition_15),
    .io_spriteYPosition_16(gameLogic_io_spriteYPosition_16),
    .io_spriteYPosition_17(gameLogic_io_spriteYPosition_17),
    .io_spriteYPosition_18(gameLogic_io_spriteYPosition_18),
    .io_spriteYPosition_19(gameLogic_io_spriteYPosition_19),
    .io_spriteYPosition_20(gameLogic_io_spriteYPosition_20),
    .io_spriteYPosition_21(gameLogic_io_spriteYPosition_21),
    .io_spriteYPosition_22(gameLogic_io_spriteYPosition_22),
    .io_spriteYPosition_23(gameLogic_io_spriteYPosition_23),
    .io_spriteYPosition_24(gameLogic_io_spriteYPosition_24),
    .io_spriteYPosition_25(gameLogic_io_spriteYPosition_25),
    .io_spriteYPosition_26(gameLogic_io_spriteYPosition_26),
    .io_spriteYPosition_27(gameLogic_io_spriteYPosition_27),
    .io_spriteYPosition_28(gameLogic_io_spriteYPosition_28),
    .io_spriteYPosition_29(gameLogic_io_spriteYPosition_29),
    .io_spriteYPosition_30(gameLogic_io_spriteYPosition_30),
    .io_spriteYPosition_31(gameLogic_io_spriteYPosition_31),
    .io_spriteYPosition_32(gameLogic_io_spriteYPosition_32),
    .io_spriteYPosition_33(gameLogic_io_spriteYPosition_33),
    .io_spriteYPosition_41(gameLogic_io_spriteYPosition_41),
    .io_spriteYPosition_42(gameLogic_io_spriteYPosition_42),
    .io_spriteYPosition_43(gameLogic_io_spriteYPosition_43),
    .io_spriteYPosition_122(gameLogic_io_spriteYPosition_122),
    .io_spriteYPosition_123(gameLogic_io_spriteYPosition_123),
    .io_spriteYPosition_124(gameLogic_io_spriteYPosition_124),
    .io_spriteYPosition_125(gameLogic_io_spriteYPosition_125),
    .io_spriteYPosition_126(gameLogic_io_spriteYPosition_126),
    .io_spriteYPosition_127(gameLogic_io_spriteYPosition_127),
    .io_spriteVisible_0(gameLogic_io_spriteVisible_0),
    .io_spriteVisible_1(gameLogic_io_spriteVisible_1),
    .io_spriteVisible_2(gameLogic_io_spriteVisible_2),
    .io_spriteVisible_3(gameLogic_io_spriteVisible_3),
    .io_spriteVisible_4(gameLogic_io_spriteVisible_4),
    .io_spriteVisible_5(gameLogic_io_spriteVisible_5),
    .io_spriteVisible_6(gameLogic_io_spriteVisible_6),
    .io_spriteVisible_7(gameLogic_io_spriteVisible_7),
    .io_spriteVisible_8(gameLogic_io_spriteVisible_8),
    .io_spriteVisible_9(gameLogic_io_spriteVisible_9),
    .io_spriteVisible_10(gameLogic_io_spriteVisible_10),
    .io_spriteVisible_11(gameLogic_io_spriteVisible_11),
    .io_spriteVisible_12(gameLogic_io_spriteVisible_12),
    .io_spriteVisible_13(gameLogic_io_spriteVisible_13),
    .io_spriteVisible_14(gameLogic_io_spriteVisible_14),
    .io_spriteVisible_15(gameLogic_io_spriteVisible_15),
    .io_spriteVisible_16(gameLogic_io_spriteVisible_16),
    .io_spriteVisible_17(gameLogic_io_spriteVisible_17),
    .io_spriteVisible_18(gameLogic_io_spriteVisible_18),
    .io_spriteVisible_19(gameLogic_io_spriteVisible_19),
    .io_spriteVisible_20(gameLogic_io_spriteVisible_20),
    .io_spriteVisible_21(gameLogic_io_spriteVisible_21),
    .io_spriteVisible_22(gameLogic_io_spriteVisible_22),
    .io_spriteVisible_23(gameLogic_io_spriteVisible_23),
    .io_spriteVisible_24(gameLogic_io_spriteVisible_24),
    .io_spriteVisible_25(gameLogic_io_spriteVisible_25),
    .io_spriteVisible_26(gameLogic_io_spriteVisible_26),
    .io_spriteVisible_27(gameLogic_io_spriteVisible_27),
    .io_spriteVisible_28(gameLogic_io_spriteVisible_28),
    .io_spriteVisible_29(gameLogic_io_spriteVisible_29),
    .io_spriteVisible_30(gameLogic_io_spriteVisible_30),
    .io_spriteVisible_31(gameLogic_io_spriteVisible_31),
    .io_spriteVisible_32(gameLogic_io_spriteVisible_32),
    .io_spriteVisible_33(gameLogic_io_spriteVisible_33),
    .io_spriteVisible_41(gameLogic_io_spriteVisible_41),
    .io_spriteVisible_42(gameLogic_io_spriteVisible_42),
    .io_spriteVisible_43(gameLogic_io_spriteVisible_43),
    .io_spriteVisible_44(gameLogic_io_spriteVisible_44),
    .io_spriteVisible_45(gameLogic_io_spriteVisible_45),
    .io_spriteVisible_46(gameLogic_io_spriteVisible_46),
    .io_spriteVisible_47(gameLogic_io_spriteVisible_47),
    .io_spriteVisible_48(gameLogic_io_spriteVisible_48),
    .io_spriteVisible_49(gameLogic_io_spriteVisible_49),
    .io_spriteVisible_50(gameLogic_io_spriteVisible_50),
    .io_spriteVisible_51(gameLogic_io_spriteVisible_51),
    .io_spriteVisible_55(gameLogic_io_spriteVisible_55),
    .io_spriteVisible_56(gameLogic_io_spriteVisible_56),
    .io_spriteVisible_57(gameLogic_io_spriteVisible_57),
    .io_spriteVisible_61(gameLogic_io_spriteVisible_61),
    .io_spriteVisible_62(gameLogic_io_spriteVisible_62),
    .io_spriteVisible_63(gameLogic_io_spriteVisible_63),
    .io_spriteVisible_64(gameLogic_io_spriteVisible_64),
    .io_spriteVisible_65(gameLogic_io_spriteVisible_65),
    .io_spriteVisible_66(gameLogic_io_spriteVisible_66),
    .io_spriteVisible_70(gameLogic_io_spriteVisible_70),
    .io_spriteVisible_71(gameLogic_io_spriteVisible_71),
    .io_spriteVisible_72(gameLogic_io_spriteVisible_72),
    .io_spriteFlipVertical_122(gameLogic_io_spriteFlipVertical_122),
    .io_spriteFlipVertical_123(gameLogic_io_spriteFlipVertical_123),
    .io_spriteFlipVertical_124(gameLogic_io_spriteFlipVertical_124),
    .io_spriteFlipVertical_125(gameLogic_io_spriteFlipVertical_125),
    .io_spriteFlipVertical_126(gameLogic_io_spriteFlipVertical_126),
    .io_spriteFlipVertical_127(gameLogic_io_spriteFlipVertical_127),
    .io_viewBoxX_0(gameLogic_io_viewBoxX_0),
    .io_backBufferWriteData(gameLogic_io_backBufferWriteData),
    .io_backBufferWriteAddress(gameLogic_io_backBufferWriteAddress),
    .io_backBufferWriteEnable(gameLogic_io_backBufferWriteEnable),
    .io_newFrame(gameLogic_io_newFrame),
    .io_frameUpdateDone(gameLogic_io_frameUpdateDone)
  );
  assign io_vgaRed = graphicEngineVGA_io_vgaRed; // @[GameTop.scala 109:13]
  assign io_vgaBlue = graphicEngineVGA_io_vgaBlue; // @[GameTop.scala 111:14]
  assign io_vgaGreen = graphicEngineVGA_io_vgaGreen; // @[GameTop.scala 110:15]
  assign io_Hsync = graphicEngineVGA_io_Hsync; // @[GameTop.scala 112:12]
  assign io_Vsync = graphicEngineVGA_io_Vsync; // @[GameTop.scala 113:12]
  assign io_soundOutput_0 = soundEngine_io_output_0; // @[GameTop.scala 67:18]
  assign io_missingFrameError = graphicEngineVGA_io_missingFrameError; // @[GameTop.scala 124:24]
  assign io_backBufferWriteError = graphicEngineVGA_io_backBufferWriteError; // @[GameTop.scala 125:27]
  assign io_viewBoxOutOfRangeError = graphicEngineVGA_io_viewBoxOutOfRangeError; // @[GameTop.scala 126:29]
  assign graphicEngineVGA_clock = clock;
  assign graphicEngineVGA_reset = _T_3 ? 1'h0 : 1'h1; // @[GameTop.scala 93:26]
  assign graphicEngineVGA_io_spriteXPosition_0 = gameLogic_io_spriteXPosition_0; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_1 = gameLogic_io_spriteXPosition_1; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_2 = gameLogic_io_spriteXPosition_2; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_3 = gameLogic_io_spriteXPosition_3; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_4 = gameLogic_io_spriteXPosition_4; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_5 = gameLogic_io_spriteXPosition_5; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_6 = gameLogic_io_spriteXPosition_6; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_7 = gameLogic_io_spriteXPosition_7; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_8 = gameLogic_io_spriteXPosition_8; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_9 = gameLogic_io_spriteXPosition_9; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_10 = gameLogic_io_spriteXPosition_10; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_11 = gameLogic_io_spriteXPosition_11; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_12 = gameLogic_io_spriteXPosition_12; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_13 = gameLogic_io_spriteXPosition_13; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_14 = gameLogic_io_spriteXPosition_14; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_15 = gameLogic_io_spriteXPosition_15; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_16 = gameLogic_io_spriteXPosition_16; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_17 = gameLogic_io_spriteXPosition_17; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_18 = gameLogic_io_spriteXPosition_18; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_19 = gameLogic_io_spriteXPosition_19; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_20 = gameLogic_io_spriteXPosition_20; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_21 = gameLogic_io_spriteXPosition_21; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_22 = gameLogic_io_spriteXPosition_22; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_23 = gameLogic_io_spriteXPosition_23; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_24 = gameLogic_io_spriteXPosition_24; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_25 = gameLogic_io_spriteXPosition_25; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_26 = gameLogic_io_spriteXPosition_26; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_27 = gameLogic_io_spriteXPosition_27; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_28 = gameLogic_io_spriteXPosition_28; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_29 = gameLogic_io_spriteXPosition_29; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_30 = gameLogic_io_spriteXPosition_30; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_31 = gameLogic_io_spriteXPosition_31; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_32 = gameLogic_io_spriteXPosition_32; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_33 = gameLogic_io_spriteXPosition_33; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_41 = gameLogic_io_spriteXPosition_41; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_42 = gameLogic_io_spriteXPosition_42; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_43 = gameLogic_io_spriteXPosition_43; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_44 = gameLogic_io_spriteXPosition_44; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_45 = gameLogic_io_spriteXPosition_45; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_46 = gameLogic_io_spriteXPosition_46; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_47 = gameLogic_io_spriteXPosition_47; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_48 = gameLogic_io_spriteXPosition_48; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_49 = gameLogic_io_spriteXPosition_49; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_50 = gameLogic_io_spriteXPosition_50; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_51 = gameLogic_io_spriteXPosition_51; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_122 = gameLogic_io_spriteXPosition_122; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_123 = gameLogic_io_spriteXPosition_123; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_124 = gameLogic_io_spriteXPosition_124; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_125 = gameLogic_io_spriteXPosition_125; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_126 = gameLogic_io_spriteXPosition_126; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteXPosition_127 = gameLogic_io_spriteXPosition_127; // @[GameTop.scala 129:39]
  assign graphicEngineVGA_io_spriteYPosition_0 = gameLogic_io_spriteYPosition_0; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_1 = gameLogic_io_spriteYPosition_1; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_2 = gameLogic_io_spriteYPosition_2; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_3 = gameLogic_io_spriteYPosition_3; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_4 = gameLogic_io_spriteYPosition_4; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_5 = gameLogic_io_spriteYPosition_5; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_6 = gameLogic_io_spriteYPosition_6; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_7 = gameLogic_io_spriteYPosition_7; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_8 = gameLogic_io_spriteYPosition_8; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_9 = gameLogic_io_spriteYPosition_9; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_10 = gameLogic_io_spriteYPosition_10; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_11 = gameLogic_io_spriteYPosition_11; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_12 = gameLogic_io_spriteYPosition_12; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_13 = gameLogic_io_spriteYPosition_13; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_14 = gameLogic_io_spriteYPosition_14; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_15 = gameLogic_io_spriteYPosition_15; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_16 = gameLogic_io_spriteYPosition_16; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_17 = gameLogic_io_spriteYPosition_17; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_18 = gameLogic_io_spriteYPosition_18; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_19 = gameLogic_io_spriteYPosition_19; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_20 = gameLogic_io_spriteYPosition_20; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_21 = gameLogic_io_spriteYPosition_21; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_22 = gameLogic_io_spriteYPosition_22; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_23 = gameLogic_io_spriteYPosition_23; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_24 = gameLogic_io_spriteYPosition_24; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_25 = gameLogic_io_spriteYPosition_25; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_26 = gameLogic_io_spriteYPosition_26; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_27 = gameLogic_io_spriteYPosition_27; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_28 = gameLogic_io_spriteYPosition_28; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_29 = gameLogic_io_spriteYPosition_29; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_30 = gameLogic_io_spriteYPosition_30; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_31 = gameLogic_io_spriteYPosition_31; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_32 = gameLogic_io_spriteYPosition_32; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_33 = gameLogic_io_spriteYPosition_33; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_41 = gameLogic_io_spriteYPosition_41; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_42 = gameLogic_io_spriteYPosition_42; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_43 = gameLogic_io_spriteYPosition_43; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_122 = gameLogic_io_spriteYPosition_122; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_123 = gameLogic_io_spriteYPosition_123; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_124 = gameLogic_io_spriteYPosition_124; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_125 = gameLogic_io_spriteYPosition_125; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_126 = gameLogic_io_spriteYPosition_126; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteYPosition_127 = gameLogic_io_spriteYPosition_127; // @[GameTop.scala 130:39]
  assign graphicEngineVGA_io_spriteVisible_0 = gameLogic_io_spriteVisible_0; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_1 = gameLogic_io_spriteVisible_1; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_2 = gameLogic_io_spriteVisible_2; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_3 = gameLogic_io_spriteVisible_3; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_4 = gameLogic_io_spriteVisible_4; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_5 = gameLogic_io_spriteVisible_5; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_6 = gameLogic_io_spriteVisible_6; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_7 = gameLogic_io_spriteVisible_7; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_8 = gameLogic_io_spriteVisible_8; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_9 = gameLogic_io_spriteVisible_9; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_10 = gameLogic_io_spriteVisible_10; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_11 = gameLogic_io_spriteVisible_11; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_12 = gameLogic_io_spriteVisible_12; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_13 = gameLogic_io_spriteVisible_13; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_14 = gameLogic_io_spriteVisible_14; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_15 = gameLogic_io_spriteVisible_15; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_16 = gameLogic_io_spriteVisible_16; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_17 = gameLogic_io_spriteVisible_17; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_18 = gameLogic_io_spriteVisible_18; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_19 = gameLogic_io_spriteVisible_19; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_20 = gameLogic_io_spriteVisible_20; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_21 = gameLogic_io_spriteVisible_21; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_22 = gameLogic_io_spriteVisible_22; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_23 = gameLogic_io_spriteVisible_23; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_24 = gameLogic_io_spriteVisible_24; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_25 = gameLogic_io_spriteVisible_25; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_26 = gameLogic_io_spriteVisible_26; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_27 = gameLogic_io_spriteVisible_27; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_28 = gameLogic_io_spriteVisible_28; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_29 = gameLogic_io_spriteVisible_29; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_30 = gameLogic_io_spriteVisible_30; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_31 = gameLogic_io_spriteVisible_31; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_32 = gameLogic_io_spriteVisible_32; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_33 = gameLogic_io_spriteVisible_33; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_41 = gameLogic_io_spriteVisible_41; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_42 = gameLogic_io_spriteVisible_42; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_43 = gameLogic_io_spriteVisible_43; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_44 = gameLogic_io_spriteVisible_44; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_45 = gameLogic_io_spriteVisible_45; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_46 = gameLogic_io_spriteVisible_46; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_47 = gameLogic_io_spriteVisible_47; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_48 = gameLogic_io_spriteVisible_48; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_49 = gameLogic_io_spriteVisible_49; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_50 = gameLogic_io_spriteVisible_50; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_51 = gameLogic_io_spriteVisible_51; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_55 = gameLogic_io_spriteVisible_55; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_56 = gameLogic_io_spriteVisible_56; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_57 = gameLogic_io_spriteVisible_57; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_61 = gameLogic_io_spriteVisible_61; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_62 = gameLogic_io_spriteVisible_62; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_63 = gameLogic_io_spriteVisible_63; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_64 = gameLogic_io_spriteVisible_64; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_65 = gameLogic_io_spriteVisible_65; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_66 = gameLogic_io_spriteVisible_66; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_70 = gameLogic_io_spriteVisible_70; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_71 = gameLogic_io_spriteVisible_71; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteVisible_72 = gameLogic_io_spriteVisible_72; // @[GameTop.scala 131:37]
  assign graphicEngineVGA_io_spriteFlipVertical_122 = gameLogic_io_spriteFlipVertical_122; // @[GameTop.scala 133:42]
  assign graphicEngineVGA_io_spriteFlipVertical_123 = gameLogic_io_spriteFlipVertical_123; // @[GameTop.scala 133:42]
  assign graphicEngineVGA_io_spriteFlipVertical_124 = gameLogic_io_spriteFlipVertical_124; // @[GameTop.scala 133:42]
  assign graphicEngineVGA_io_spriteFlipVertical_125 = gameLogic_io_spriteFlipVertical_125; // @[GameTop.scala 133:42]
  assign graphicEngineVGA_io_spriteFlipVertical_126 = gameLogic_io_spriteFlipVertical_126; // @[GameTop.scala 133:42]
  assign graphicEngineVGA_io_spriteFlipVertical_127 = gameLogic_io_spriteFlipVertical_127; // @[GameTop.scala 133:42]
  assign graphicEngineVGA_io_viewBoxX_0 = gameLogic_io_viewBoxX_0; // @[GameTop.scala 136:32]
  assign graphicEngineVGA_io_backBufferWriteData = gameLogic_io_backBufferWriteData; // @[GameTop.scala 140:43]
  assign graphicEngineVGA_io_backBufferWriteAddress = gameLogic_io_backBufferWriteAddress; // @[GameTop.scala 141:46]
  assign graphicEngineVGA_io_backBufferWriteEnable = gameLogic_io_backBufferWriteEnable; // @[GameTop.scala 142:45]
  assign graphicEngineVGA_io_frameUpdateDone = gameLogic_io_frameUpdateDone; // @[GameTop.scala 146:39]
  assign soundEngine_clock = clock;
  assign soundEngine_reset = reset;
  assign soundEngine_io_input = gameLogic_io_songInput; // @[GameTop.scala 64:24]
  assign gameLogic_clock = clock;
  assign gameLogic_reset = _T_3 ? 1'h0 : 1'h1; // @[GameTop.scala 94:19]
  assign gameLogic_io_btnC = btnCState; // @[GameTop.scala 102:21]
  assign gameLogic_io_btnU = btnUState; // @[GameTop.scala 103:21]
  assign gameLogic_io_btnL = btnLState; // @[GameTop.scala 104:21]
  assign gameLogic_io_btnR = btnRState; // @[GameTop.scala 105:21]
  assign gameLogic_io_btnD = btnDState; // @[GameTop.scala 106:21]
  assign gameLogic_io_sw_0 = _T_18; // @[GameTop.scala 117:24]
  assign gameLogic_io_sw_1 = _T_21; // @[GameTop.scala 117:24]
  assign gameLogic_io_sw_2 = _T_24; // @[GameTop.scala 117:24]
  assign gameLogic_io_sw_7 = _T_39; // @[GameTop.scala 117:24]
  assign gameLogic_io_newFrame = graphicEngineVGA_io_newFrame; // @[GameTop.scala 145:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounceCounter = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  resetReleaseCounter = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  _T_7_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_7_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_7_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btnCState = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_9_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_9_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_9_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btnUState = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_11_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_11_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_11_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btnLState = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_13_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_13_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_13_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btnRState = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_15_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_15_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_15_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  btnDState = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_17_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_17_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_17_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_18 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_20_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_20_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_20_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_21 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_23_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_23_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_23_2 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_24 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_38_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_38_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_38_2 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_39 = _RAND_37[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      debounceCounter <= 21'h0;
    end else if (debounceSampleEn) begin
      debounceCounter <= 21'h0;
    end else begin
      debounceCounter <= _T_2;
    end
    if (reset) begin
      resetReleaseCounter <= 22'h0;
    end else if (!(_T_3)) begin
      resetReleaseCounter <= _T_5;
    end
    if (reset) begin
      _T_7_0 <= 1'h0;
    end else begin
      _T_7_0 <= _T_7_1;
    end
    if (reset) begin
      _T_7_1 <= 1'h0;
    end else begin
      _T_7_1 <= _T_7_2;
    end
    if (reset) begin
      _T_7_2 <= 1'h0;
    end else begin
      _T_7_2 <= io_btnC;
    end
    if (reset) begin
      btnCState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnCState <= _T_7_0;
    end
    if (reset) begin
      _T_9_0 <= 1'h0;
    end else begin
      _T_9_0 <= _T_9_1;
    end
    if (reset) begin
      _T_9_1 <= 1'h0;
    end else begin
      _T_9_1 <= _T_9_2;
    end
    if (reset) begin
      _T_9_2 <= 1'h0;
    end else begin
      _T_9_2 <= io_btnU;
    end
    if (reset) begin
      btnUState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnUState <= _T_9_0;
    end
    if (reset) begin
      _T_11_0 <= 1'h0;
    end else begin
      _T_11_0 <= _T_11_1;
    end
    if (reset) begin
      _T_11_1 <= 1'h0;
    end else begin
      _T_11_1 <= _T_11_2;
    end
    if (reset) begin
      _T_11_2 <= 1'h0;
    end else begin
      _T_11_2 <= io_btnL;
    end
    if (reset) begin
      btnLState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnLState <= _T_11_0;
    end
    if (reset) begin
      _T_13_0 <= 1'h0;
    end else begin
      _T_13_0 <= _T_13_1;
    end
    if (reset) begin
      _T_13_1 <= 1'h0;
    end else begin
      _T_13_1 <= _T_13_2;
    end
    if (reset) begin
      _T_13_2 <= 1'h0;
    end else begin
      _T_13_2 <= io_btnR;
    end
    if (reset) begin
      btnRState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnRState <= _T_13_0;
    end
    if (reset) begin
      _T_15_0 <= 1'h0;
    end else begin
      _T_15_0 <= _T_15_1;
    end
    if (reset) begin
      _T_15_1 <= 1'h0;
    end else begin
      _T_15_1 <= _T_15_2;
    end
    if (reset) begin
      _T_15_2 <= 1'h0;
    end else begin
      _T_15_2 <= io_btnD;
    end
    if (reset) begin
      btnDState <= 1'h0;
    end else if (debounceSampleEn) begin
      btnDState <= _T_15_0;
    end
    if (reset) begin
      _T_17_0 <= 1'h0;
    end else begin
      _T_17_0 <= _T_17_1;
    end
    if (reset) begin
      _T_17_1 <= 1'h0;
    end else begin
      _T_17_1 <= _T_17_2;
    end
    if (reset) begin
      _T_17_2 <= 1'h0;
    end else begin
      _T_17_2 <= io_sw_0;
    end
    if (reset) begin
      _T_18 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_18 <= _T_17_0;
    end
    if (reset) begin
      _T_20_0 <= 1'h0;
    end else begin
      _T_20_0 <= _T_20_1;
    end
    if (reset) begin
      _T_20_1 <= 1'h0;
    end else begin
      _T_20_1 <= _T_20_2;
    end
    if (reset) begin
      _T_20_2 <= 1'h0;
    end else begin
      _T_20_2 <= io_sw_1;
    end
    if (reset) begin
      _T_21 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_21 <= _T_20_0;
    end
    if (reset) begin
      _T_23_0 <= 1'h0;
    end else begin
      _T_23_0 <= _T_23_1;
    end
    if (reset) begin
      _T_23_1 <= 1'h0;
    end else begin
      _T_23_1 <= _T_23_2;
    end
    if (reset) begin
      _T_23_2 <= 1'h0;
    end else begin
      _T_23_2 <= io_sw_2;
    end
    if (reset) begin
      _T_24 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_24 <= _T_23_0;
    end
    if (reset) begin
      _T_38_0 <= 1'h0;
    end else begin
      _T_38_0 <= _T_38_1;
    end
    if (reset) begin
      _T_38_1 <= 1'h0;
    end else begin
      _T_38_1 <= _T_38_2;
    end
    if (reset) begin
      _T_38_2 <= 1'h0;
    end else begin
      _T_38_2 <= io_sw_7;
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else if (debounceSampleEn) begin
      _T_39 <= _T_38_0;
    end
  end
endmodule
module Top(
  input        clock,
  input        reset,
  input        io_btnC,
  input        io_btnU,
  input        io_btnL,
  input        io_btnR,
  input        io_btnD,
  output [3:0] io_vgaRed,
  output [3:0] io_vgaGreen,
  output [3:0] io_vgaBlue,
  output       io_Hsync,
  output       io_Vsync,
  input        io_sw_0,
  input        io_sw_1,
  input        io_sw_2,
  input        io_sw_3,
  input        io_sw_4,
  input        io_sw_5,
  input        io_sw_6,
  input        io_sw_7,
  output       io_led_0,
  output       io_led_1,
  output       io_led_2,
  output       io_led_3,
  output       io_led_4,
  output       io_led_5,
  output       io_led_6,
  output       io_led_7,
  output       io_soundOutput_0,
  output       io_missingFrameError,
  output       io_backBufferWriteError,
  output       io_viewBoxOutOfRangeError
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  gameTop_clock; // @[Top.scala 42:23]
  wire  gameTop_reset; // @[Top.scala 42:23]
  wire  gameTop_io_btnC; // @[Top.scala 42:23]
  wire  gameTop_io_btnU; // @[Top.scala 42:23]
  wire  gameTop_io_btnL; // @[Top.scala 42:23]
  wire  gameTop_io_btnR; // @[Top.scala 42:23]
  wire  gameTop_io_btnD; // @[Top.scala 42:23]
  wire [3:0] gameTop_io_vgaRed; // @[Top.scala 42:23]
  wire [3:0] gameTop_io_vgaBlue; // @[Top.scala 42:23]
  wire [3:0] gameTop_io_vgaGreen; // @[Top.scala 42:23]
  wire  gameTop_io_Hsync; // @[Top.scala 42:23]
  wire  gameTop_io_Vsync; // @[Top.scala 42:23]
  wire  gameTop_io_sw_0; // @[Top.scala 42:23]
  wire  gameTop_io_sw_1; // @[Top.scala 42:23]
  wire  gameTop_io_sw_2; // @[Top.scala 42:23]
  wire  gameTop_io_sw_7; // @[Top.scala 42:23]
  wire  gameTop_io_soundOutput_0; // @[Top.scala 42:23]
  wire  gameTop_io_missingFrameError; // @[Top.scala 42:23]
  wire  gameTop_io_backBufferWriteError; // @[Top.scala 42:23]
  wire  gameTop_io_viewBoxOutOfRangeError; // @[Top.scala 42:23]
  reg  _T_1; // @[Top.scala 47:48]
  reg  _T_2; // @[Top.scala 47:40]
  reg  _T_3; // @[Top.scala 47:32]
  reg  pipeResetReg_0; // @[Top.scala 52:25]
  reg  pipeResetReg_1; // @[Top.scala 52:25]
  reg  pipeResetReg_2; // @[Top.scala 52:25]
  reg  pipeResetReg_3; // @[Top.scala 52:25]
  reg  pipeResetReg_4; // @[Top.scala 52:25]
  wire [4:0] _T_7 = {pipeResetReg_4,pipeResetReg_3,pipeResetReg_2,pipeResetReg_1,pipeResetReg_0}; // @[Top.scala 57:33]
  GameTop gameTop ( // @[Top.scala 42:23]
    .clock(gameTop_clock),
    .reset(gameTop_reset),
    .io_btnC(gameTop_io_btnC),
    .io_btnU(gameTop_io_btnU),
    .io_btnL(gameTop_io_btnL),
    .io_btnR(gameTop_io_btnR),
    .io_btnD(gameTop_io_btnD),
    .io_vgaRed(gameTop_io_vgaRed),
    .io_vgaBlue(gameTop_io_vgaBlue),
    .io_vgaGreen(gameTop_io_vgaGreen),
    .io_Hsync(gameTop_io_Hsync),
    .io_Vsync(gameTop_io_Vsync),
    .io_sw_0(gameTop_io_sw_0),
    .io_sw_1(gameTop_io_sw_1),
    .io_sw_2(gameTop_io_sw_2),
    .io_sw_7(gameTop_io_sw_7),
    .io_soundOutput_0(gameTop_io_soundOutput_0),
    .io_missingFrameError(gameTop_io_missingFrameError),
    .io_backBufferWriteError(gameTop_io_backBufferWriteError),
    .io_viewBoxOutOfRangeError(gameTop_io_viewBoxOutOfRangeError)
  );
  assign io_vgaRed = gameTop_io_vgaRed; // @[Top.scala 60:14]
  assign io_vgaGreen = gameTop_io_vgaGreen; // @[Top.scala 60:14]
  assign io_vgaBlue = gameTop_io_vgaBlue; // @[Top.scala 60:14]
  assign io_Hsync = gameTop_io_Hsync; // @[Top.scala 60:14]
  assign io_Vsync = gameTop_io_Vsync; // @[Top.scala 60:14]
  assign io_led_0 = 1'h0; // @[Top.scala 60:14]
  assign io_led_1 = 1'h0; // @[Top.scala 60:14]
  assign io_led_2 = 1'h0; // @[Top.scala 60:14]
  assign io_led_3 = 1'h0; // @[Top.scala 60:14]
  assign io_led_4 = 1'h0; // @[Top.scala 60:14]
  assign io_led_5 = 1'h0; // @[Top.scala 60:14]
  assign io_led_6 = 1'h0; // @[Top.scala 60:14]
  assign io_led_7 = 1'h0; // @[Top.scala 60:14]
  assign io_soundOutput_0 = gameTop_io_soundOutput_0; // @[Top.scala 60:14]
  assign io_missingFrameError = gameTop_io_missingFrameError; // @[Top.scala 60:14]
  assign io_backBufferWriteError = gameTop_io_backBufferWriteError; // @[Top.scala 60:14]
  assign io_viewBoxOutOfRangeError = gameTop_io_viewBoxOutOfRangeError; // @[Top.scala 60:14]
  assign gameTop_clock = clock;
  assign gameTop_reset = |_T_7; // @[Top.scala 57:17]
  assign gameTop_io_btnC = io_btnC; // @[Top.scala 60:14]
  assign gameTop_io_btnU = io_btnU; // @[Top.scala 60:14]
  assign gameTop_io_btnL = io_btnL; // @[Top.scala 60:14]
  assign gameTop_io_btnR = io_btnR; // @[Top.scala 60:14]
  assign gameTop_io_btnD = io_btnD; // @[Top.scala 60:14]
  assign gameTop_io_sw_0 = io_sw_0; // @[Top.scala 60:14]
  assign gameTop_io_sw_1 = io_sw_1; // @[Top.scala 60:14]
  assign gameTop_io_sw_2 = io_sw_2; // @[Top.scala 60:14]
  assign gameTop_io_sw_7 = io_sw_7; // @[Top.scala 60:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_2 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pipeResetReg_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pipeResetReg_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pipeResetReg_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pipeResetReg_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pipeResetReg_4 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= reset;
    _T_2 <= _T_1;
    _T_3 <= _T_2;
    pipeResetReg_0 <= pipeResetReg_1;
    pipeResetReg_1 <= pipeResetReg_2;
    pipeResetReg_2 <= pipeResetReg_3;
    pipeResetReg_3 <= pipeResetReg_4;
    pipeResetReg_4 <= ~_T_3;
  end
endmodule
